library ieee;
use ieee.std_logic_1164.all;

entity reference is
   port (
      clear    : in  bit;
      start    : in  bit;
      y0       : in  bit;
      y1       : in  bit;
      y2       : in  bit;
      y3       : in  bit;
      senddata : out bit_vector (3 downto 0);
      match    : out bit_vector (3 downto 0)
      );
end reference;

architecture verify of reference is

type senddata_rom is array (000 to 2499) of bit_vector (3 downto 0);
constant senddata_tbl : senddata_rom :=
(

 B"0010", B"0001", B"1101", B"1011", 
 B"1000", B"1011", B"1101", B"1100", 
 B"0010", B"0011", B"1100", B"1010", 
 B"1001", B"1111", B"0110", B"0010", 
 B"1100", B"1000", B"0001", B"1010", 
 B"0110", B"1011", B"0101", B"0001", 
 B"1100", B"1001", B"1100", B"1000", 
 B"0110", B"1101", B"0000", B"0100", 
 B"0000", B"0110", B"1101", B"1011", 
 B"0000", B"1001", B"1001", B"1000", 
 B"0110", B"1100", B"0110", B"1101", 
 B"1101", B"1011", B"0101", B"1101", 
 B"1111", B"0110", B"1000", B"0010", 
 B"1111", B"0110", B"0000", B"1110", 
 B"0001", B"0101", B"0111", B"1111", 
 B"0100", B"1010", B"1011", B"0111", 
 B"0011", B"1101", B"1000", B"1000", 
 B"0001", B"1000", B"1110", B"0110", 
 B"1111", B"1101", B"0000", B"0000", 
 B"1111", B"1010", B"1001", B"0011", 
 B"1110", B"0010", B"0010", B"0011", 
 B"1000", B"1101", B"1101", B"0000", 
 B"0000", B"1001", B"1010", B"1010", 
 B"0000", B"0111", B"0001", B"1111", 
 B"1010", B"0110", B"0100", B"0000", 
 B"1011", B"1100", B"0000", B"0011", 
 B"1111", B"0001", B"0000", B"0000", 
 B"1011", B"0100", B"1101", B"0011", 
 B"0001", B"1000", B"0101", B"0000", 
 B"0100", B"1111", B"0100", B"0010", 
 B"0101", B"0000", B"0001", B"0100", 
 B"1000", B"0000", B"1101", B"1100", 
 B"1110", B"1100", B"1001", B"0010", 
 B"0101", B"0001", B"0101", B"1001", 
 B"0011", B"1010", B"0111", B"1101", 
 B"0010", B"1111", B"1010", B"0011", 
 B"0011", B"0010", B"0111", B"0010", 
 B"0000", B"0001", B"0110", B"1100", 
 B"0001", B"0110", B"1110", B"0110", 
 B"1101", B"0001", B"1101", B"0001", 
 B"0011", B"1000", B"1001", B"1010", 
 B"0110", B"1101", B"0110", B"1010", 
 B"0011", B"0010", B"1110", B"1101", 
 B"1011", B"0010", B"1110", B"1000", 
 B"0010", B"1111", B"0010", B"0110", 
 B"1110", B"1100", B"0000", B"0000", 
 B"0000", B"0110", B"1110", B"0101", 
 B"1010", B"1000", B"0100", B"0001", 
 B"0101", B"0110", B"1101", B"1011", 
 B"1000", B"1111", B"1111", B"1101", 
 B"0001", B"1011", B"1000", B"0011", 
 B"0010", B"0100", B"0010", B"0010", 
 B"0010", B"0101", B"0111", B"1101", 
 B"1000", B"1101", B"1001", B"1001", 
 B"0101", B"0011", B"0100", B"0000", 
 B"1100", B"1100", B"1000", B"1001", 
 B"0000", B"1110", B"0110", B"1101", 
 B"0010", B"0000", B"1111", B"1010", 
 B"1010", B"0100", B"1101", B"0010", 
 B"1001", B"1001", B"1011", B"1000", 
 B"0000", B"1001", B"1110", B"0000", 
 B"0110", B"1000", B"0101", B"0010", 
 B"1100", B"0100", B"1000", B"0110", 
 B"0100", B"1111", B"0011", B"0101", 
 B"0000", B"1100", B"0110", B"1110", 
 B"1111", B"1000", B"1000", B"0110", 
 B"1000", B"1000", B"1100", B"1000", 
 B"1100", B"0011", B"0110", B"1001", 
 B"0101", B"0011", B"0111", B"0100", 
 B"0010", B"1011", B"1001", B"0111", 
 B"1110", B"0001", B"1001", B"0110", 
 B"1001", B"0111", B"1111", B"0010", 
 B"1010", B"0011", B"0101", B"1010", 
 B"0000", B"0000", B"0001", B"0110", 
 B"1111", B"0010", B"0100", B"1100", 
 B"0100", B"0001", B"0000", B"1010", 
 B"1001", B"1011", B"0101", B"1101", 
 B"1100", B"1010", B"0010", B"1101", 
 B"1111", B"1000", B"0111", B"0101", 
 B"0010", B"1101", B"0111", B"1110", 
 B"1011", B"0110", B"0101", B"1010", 
 B"1001", B"0001", B"0001", B"1000", 
 B"0100", B"1010", B"1111", B"1100", 
 B"1000", B"0101", B"1010", B"0011", 
 B"0010", B"1010", B"1010", B"0110", 
 B"0101", B"0000", B"0011", B"0011", 
 B"0110", B"0011", B"1100", B"1111", 
 B"0001", B"1101", B"1011", B"1111", 
 B"1100", B"1000", B"0010", B"1100", 
 B"0010", B"1100", B"0001", B"1101", 
 B"0111", B"0001", B"1110", B"1010", 
 B"0010", B"1111", B"0101", B"1011", 
 B"1110", B"0001", B"0001", B"1000", 
 B"1000", B"1000", B"1011", B"0101", 
 B"1000", B"1011", B"0011", B"0001", 
 B"1110", B"1111", B"0111", B"0010", 
 B"0101", B"0110", B"0000", B"1110", 
 B"0000", B"0110", B"1011", B"0101", 
 B"0001", B"0001", B"1111", B"1100", 
 B"1110", B"0000", B"0101", B"1011", 
 B"1011", B"0000", B"0110", B"0111", 
 B"0111", B"1110", B"0011", B"0000", 
 B"1100", B"0110", B"0000", B"1000", 
 B"0010", B"0100", B"1101", B"0000", 
 B"0000", B"0001", B"0100", B"1101", 
 B"0011", B"1001", B"0110", B"1001", 
 B"0000", B"0000", B"0001", B"1011", 
 B"1000", B"1001", B"0000", B"1000", 
 B"1101", B"0111", B"0110", B"0100", 
 B"1011", B"0010", B"0000", B"0100", 
 B"1010", B"1101", B"1011", B"1100", 
 B"0111", B"1111", B"0110", B"0011", 
 B"0001", B"0100", B"0001", B"1010", 
 B"1011", B"0110", B"1111", B"1010", 
 B"1110", B"0010", B"1000", B"0100", 
 B"0010", B"1010", B"1010", B"1010", 
 B"0001", B"1010", B"0000", B"1010", 
 B"0101", B"1011", B"0000", B"0100", 
 B"1000", B"1111", B"0100", B"1010", 
 B"1111", B"1000", B"1110", B"0111", 
 B"1110", B"1011", B"0000", B"1100", 
 B"0011", B"0000", B"1011", B"1100", 
 B"0010", B"1000", B"1011", B"0110", 
 B"1000", B"1111", B"1000", B"0110", 
 B"1100", B"1001", B"1101", B"1001", 
 B"0010", B"0100", B"0101", B"0101", 
 B"1010", B"0000", B"1000", B"1010", 
 B"1100", B"0110", B"0110", B"1100", 
 B"0011", B"0010", B"0000", B"0100", 
 B"0010", B"1010", B"1010", B"0101", 
 B"0110", B"1000", B"0001", B"0100", 
 B"1111", B"0011", B"0111", B"1001", 
 B"0111", B"0110", B"1100", B"1010", 
 B"1001", B"0011", B"0000", B"0010", 
 B"0110", B"0000", B"1100", B"1101", 
 B"0100", B"0010", B"1110", B"0011", 
 B"0001", B"1011", B"0000", B"1010", 
 B"0011", B"0011", B"0111", B"0100", 
 B"0001", B"1100", B"1000", B"1101", 
 B"0100", B"1101", B"0010", B"1011", 
 B"1010", B"1011", B"0011", B"1000", 
 B"1000", B"0010", B"1010", B"0010", 
 B"0110", B"1100", B"1110", B"0010", 
 B"0110", B"0001", B"0111", B"1101", 
 B"1101", B"1111", B"0010", B"0001", 
 B"0011", B"0110", B"0100", B"0101", 
 B"1001", B"0011", B"0000", B"0101", 
 B"1111", B"0010", B"1110", B"1010", 
 B"1111", B"0011", B"1101", B"0011", 
 B"0000", B"0101", B"0011", B"0100", 
 B"0101", B"0111", B"1100", B"0101", 
 B"0010", B"1101", B"0010", B"1100", 
 B"1110", B"1110", B"0011", B"0101", 
 B"1001", B"0111", B"0001", B"0011", 
 B"1000", B"0010", B"0001", B"1000", 
 B"1010", B"0110", B"0101", B"0010", 
 B"0101", B"0010", B"1011", B"1111", 
 B"1110", B"0100", B"0110", B"1001", 
 B"0110", B"0111", B"0111", B"1000", 
 B"0001", B"0111", B"1101", B"1110", 
 B"1011", B"1111", B"0010", B"0100", 
 B"1110", B"0111", B"0000", B"1011", 
 B"0001", B"0010", B"0000", B"1011", 
 B"0000", B"0101", B"0001", B"1111", 
 B"0000", B"1101", B"1101", B"0010", 
 B"1011", B"1110", B"1110", B"0001", 
 B"0010", B"1011", B"0011", B"1101", 
 B"0101", B"1011", B"1100", B"1100", 
 B"1001", B"0101", B"0000", B"0111", 
 B"1111", B"1000", B"0010", B"0100", 
 B"1100", B"1001", B"0111", B"1001", 
 B"0101", B"0000", B"1110", B"1000", 
 B"1011", B"0111", B"0101", B"1001", 
 B"0101", B"0000", B"1100", B"0111", 
 B"1001", B"1110", B"1001", B"1011", 
 B"1010", B"0011", B"1101", B"1101", 
 B"0101", B"0101", B"1110", B"1011", 
 B"1011", B"1101", B"0111", B"0101", 
 B"1010", B"1101", B"1101", B"1000", 
 B"1101", B"0001", B"1110", B"0101", 
 B"0100", B"0001", B"0010", B"1011", 
 B"1001", B"1001", B"1110", B"1101", 
 B"0101", B"0110", B"0001", B"1101", 
 B"0011", B"0111", B"0110", B"0001", 
 B"0011", B"1111", B"0101", B"1101", 
 B"1111", B"0000", B"1000", B"1001", 
 B"1111", B"1100", B"0110", B"0001", 
 B"1100", B"1010", B"1111", B"0011", 
 B"1000", B"0100", B"1101", B"0100", 
 B"0100", B"0111", B"1011", B"1110", 
 B"0101", B"0101", B"1011", B"1001", 
 B"0001", B"0110", B"0110", B"1111", 
 B"1110", B"1100", B"1100", B"1011", 
 B"1000", B"1010", B"1100", B"1001", 
 B"0101", B"0010", B"0010", B"0011", 
 B"1001", B"0010", B"0010", B"0111", 
 B"1111", B"0100", B"0001", B"0000", 
 B"1001", B"1100", B"0010", B"1010", 
 B"0100", B"0110", B"0010", B"0001", 
 B"1111", B"0100", B"0001", B"0101", 
 B"0001", B"0010", B"0111", B"0010", 
 B"1110", B"0100", B"0001", B"1100", 
 B"0111", B"1100", B"1010", B"0011", 
 B"1010", B"1110", B"0100", B"0101", 
 B"0001", B"0000", B"0100", B"1000", 
 B"1001", B"0010", B"0100", B"0000", 
 B"0011", B"1111", B"1010", B"0010", 
 B"0110", B"0111", B"1110", B"0101", 
 B"1111", B"0110", B"0010", B"0011", 
 B"1101", B"0001", B"1000", B"1101", 
 B"0001", B"1111", B"1110", B"1111", 
 B"1011", B"1100", B"0001", B"0001", 
 B"1111", B"0000", B"1000", B"0000", 
 B"1111", B"1110", B"0011", B"0110", 
 B"1000", B"0101", B"0100", B"1000", 
 B"0001", B"0001", B"1001", B"0100", 
 B"1000", B"1101", B"1100", B"0000", 
 B"1101", B"1111", B"1011", B"1011", 
 B"1110", B"1100", B"0010", B"0111", 
 B"0000", B"0000", B"1101", B"1101", 
 B"0010", B"0000", B"1000", B"0100", 
 B"1001", B"1001", B"1111", B"1001", 
 B"0001", B"1110", B"1110", B"1111", 
 B"0111", B"1010", B"0000", B"1100", 
 B"0111", B"1110", B"1010", B"0100", 
 B"0100", B"0010", B"1101", B"0000", 
 B"1100", B"0011", B"1100", B"0011", 
 B"0010", B"1001", B"0010", B"1011", 
 B"0110", B"1010", B"1011", B"1110", 
 B"0001", B"0110", B"1001", B"0000", 
 B"1111", B"0100", B"0100", B"0011", 
 B"1101", B"0110", B"1101", B"0101", 
 B"0001", B"1100", B"1101", B"0100", 
 B"0001", B"1110", B"0011", B"1101", 
 B"1101", B"0000", B"1110", B"0010", 
 B"1001", B"0110", B"1000", B"0000", 
 B"1000", B"1010", B"1011", B"1000", 
 B"0110", B"0010", B"1010", B"1111", 
 B"1000", B"0011", B"1010", B"0000", 
 B"0010", B"1011", B"1110", B"1000", 
 B"0011", B"0100", B"0101", B"1001", 
 B"0100", B"0111", B"1110", B"0111", 
 B"0011", B"0111", B"0100", B"1100", 
 B"1010", B"0110", B"1011", B"1111", 
 B"1110", B"1011", B"0111", B"1110", 
 B"0011", B"0011", B"0011", B"0001", 
 B"0110", B"1110", B"1000", B"0000", 
 B"1100", B"0001", B"0100", B"0001", 
 B"0010", B"1001", B"0011", B"0100", 
 B"0011", B"0011", B"0111", B"1001", 
 B"1111", B"1101", B"0000", B"0000", 
 B"1010", B"0000", B"0110", B"0110", 
 B"0001", B"1100", B"1111", B"1100", 
 B"0000", B"1001", B"1101", B"0001", 
 B"1001", B"0101", B"0101", B"0101", 
 B"1000", B"0101", B"0001", B"1100", 
 B"1111", B"1111", B"1000", B"1110", 
 B"1000", B"0101", B"0011", B"1111", 
 B"0110", B"1001", B"1010", B"0011", 
 B"1101", B"1011", B"0010", B"1100", 
 B"0000", B"0101", B"0000", B"0011", 
 B"1110", B"1001", B"0111", B"0110", 
 B"0110", B"0011", B"1010", B"0000", 
 B"1000", B"0111", B"0111", B"1101", 
 B"1001", B"0001", B"1011", B"1100", 
 B"1101", B"0110", B"1101", B"0010", 
 B"1010", B"0001", B"0001", B"0111", 
 B"0001", B"1011", B"1100", B"1101", 
 B"0010", B"0001", B"0110", B"1101", 
 B"1111", B"0001", B"0011", B"0001", 
 B"1010", B"0100", B"0001", B"1111", 
 B"0011", B"1010", B"1011", B"1000", 
 B"1101", B"0011", B"0010", B"0001", 
 B"1110", B"0101", B"1111", B"0101", 
 B"1000", B"1001", B"0101", B"1011", 
 B"0111", B"1111", B"0001", B"0100", 
 B"1111", B"1000", B"1000", B"0111", 
 B"0101", B"0011", B"0001", B"0000", 
 B"0101", B"1101", B"1110", B"0001", 
 B"0110", B"1011", B"0110", B"0000", 
 B"1100", B"0001", B"1100", B"1101", 
 B"1111", B"0111", B"0001", B"0100", 
 B"0100", B"1100", B"1100", B"1101", 
 B"1010", B"1011", B"1010", B"1011", 
 B"1101", B"0100", B"0100", B"0011", 
 B"1111", B"1010", B"0110", B"1001", 
 B"1111", B"0110", B"0110", B"0000", 
 B"1010", B"0111", B"0111", B"0011", 
 B"0101", B"1001", B"0000", B"0111", 
 B"0110", B"1100", B"0001", B"1100", 
 B"1010", B"0101", B"0000", B"0010", 
 B"1111", B"0011", B"1001", B"1000", 
 B"0101", B"0110", B"1001", B"1110", 
 B"0111", B"1011", B"1000", B"0001", 
 B"1001", B"1110", B"1011", B"0101", 
 B"0001", B"1111", B"1111", B"0010", 
 B"1101", B"0010", B"0010", B"0001", 
 B"0100", B"0100", B"1101", B"1001", 
 B"1001", B"1100", B"1000", B"1001", 
 B"0010", B"0111", B"1010", B"0011", 
 B"0010", B"1011", B"0011", B"0110", 
 B"1010", B"0111", B"0010", B"0111", 
 B"0011", B"0011", B"0100", B"1110", 
 B"1110", B"1100", B"0001", B"0011", 
 B"0000", B"1010", B"1110", B"0010", 
 B"1001", B"1000", B"1100", B"1000", 
 B"0010", B"0001", B"0110", B"0100", 
 B"1011", B"1000", B"1111", B"1001", 
 B"0001", B"1101", B"0001", B"0000", 
 B"0101", B"0111", B"1001", B"1011", 
 B"1000", B"0111", B"1001", B"1000", 
 B"0011", B"1100", B"1000", B"1111", 
 B"1010", B"0111", B"0001", B"0101", 
 B"1001", B"1111", B"1101", B"1010", 
 B"0100", B"0010", B"0101", B"1010", 
 B"1011", B"0100", B"1000", B"0110", 
 B"1001", B"1100", B"1000", B"1100", 
 B"0011", B"1001", B"0011", B"1101", 
 B"1100", B"0000", B"1010", B"1000", 
 B"1001", B"0111", B"1001", B"1100", 
 B"0000", B"0101", B"0101", B"0010", 
 B"1011", B"0101", B"1100", B"0101", 
 B"1001", B"1010", B"1000", B"1100", 
 B"1000", B"1101", B"1101", B"0001", 
 B"0110", B"0110", B"1011", B"1010", 
 B"0010", B"1100", B"0111", B"0010", 
 B"0110", B"0001", B"0010", B"1111", 
 B"0110", B"0101", B"1111", B"0011", 
 B"1110", B"0000", B"1010", B"0110", 
 B"1101", B"0011", B"1010", B"0111", 
 B"0000", B"0110", B"0010", B"0001", 
 B"0100", B"1011", B"0011", B"0111", 
 B"0100", B"1010", B"0111", B"1110", 
 B"1100", B"1110", B"1101", B"0011", 
 B"0111", B"0010", B"0000", B"1111", 
 B"0010", B"1100", B"0110", B"0110", 
 B"0000", B"0000", B"1010", B"1101", 
 B"0100", B"0111", B"0001", B"1010", 
 B"0000", B"0011", B"1011", B"1010", 
 B"1100", B"1000", B"0101", B"1110", 
 B"1101", B"1001", B"1110", B"1111", 
 B"1110", B"0111", B"1101", B"1010", 
 B"1001", B"1010", B"1111", B"0111", 
 B"0110", B"1000", B"1010", B"0101", 
 B"1110", B"1010", B"0000", B"0111", 
 B"0110", B"1111", B"1000", B"1001", 
 B"0110", B"0101", B"0010", B"1011", 
 B"1111", B"0000", B"1100", B"0101", 
 B"0101", B"1101", B"0111", B"0111", 
 B"0101", B"0011", B"0101", B"0011", 
 B"0011", B"1000", B"1101", B"1011", 
 B"1000", B"0111", B"1010", B"1100", 
 B"1110", B"0100", B"0011", B"1110", 
 B"1001", B"1011", B"0100", B"1010", 
 B"1010", B"0101", B"1011", B"0101", 
 B"1011", B"0100", B"0110", B"0110", 
 B"1000", B"0010", B"1111", B"0010", 
 B"1111", B"1011", B"1000", B"0000", 
 B"0100", B"0110", B"0001", B"0010", 
 B"0001", B"0110", B"0100", B"1111", 
 B"0110", B"0001", B"0010", B"1001", 
 B"0011", B"0011", B"0100", B"0111", 
 B"0100", B"1111", B"0100", B"0101", 
 B"0100", B"1000", B"0011", B"1000", 
 B"0011", B"0110", B"1001", B"0101", 
 B"1001", B"1100", B"1011", B"0010", 
 B"0000", B"0010", B"0010", B"1110", 
 B"0100", B"0010", B"0100", B"0110", 
 B"1001", B"1101", B"1010", B"1111", 
 B"1101", B"0110", B"0100", B"0111", 
 B"0111", B"1000", B"0111", B"1000", 
 B"0010", B"0110", B"1000", B"1001", 
 B"0011", B"1100", B"0010", B"0010", 
 B"1111", B"0011", B"0000", B"1111", 
 B"1100", B"0001", B"1000", B"0001", 
 B"1000", B"0110", B"1010", B"1111", 
 B"0100", B"0111", B"0010", B"0111", 
 B"1001", B"0100", B"0001", B"1000", 
 B"0100", B"1110", B"0010", B"1110", 
 B"0110", B"1000", B"0110", B"0111", 
 B"0110", B"0001", B"0110", B"0001", 
 B"1101", B"1000", B"1111", B"1001", 
 B"0011", B"0011", B"1011", B"1111", 
 B"1100", B"1001", B"1101", B"1111", 
 B"0010", B"1101", B"0010", B"1010", 
 B"0100", B"1000", B"0000", B"0000", 
 B"1100", B"1011", B"0100", B"0011", 
 B"0100", B"1001", B"1001", B"0011", 
 B"1001", B"0110", B"1111", B"1011", 
 B"0001", B"1011", B"0000", B"0110", 
 B"0101", B"0111", B"0101", B"1101", 
 B"0011", B"0110", B"1100", B"1001", 
 B"1110", B"1111", B"1101", B"0110", 
 B"1010", B"0101", B"1000", B"1010", 
 B"0000", B"1011", B"1100", B"1000", 
 B"1111", B"0101", B"0111", B"1011", 
 B"0101", B"1101", B"1110", B"0101", 
 B"1000", B"0011", B"1101", B"1110", 
 B"0110", B"1100", B"1110", B"0000", 
 B"1011", B"1011", B"0000", B"0001", 
 B"0011", B"1101", B"0011", B"1111", 
 B"1000", B"1101", B"1001", B"1110", 
 B"1100", B"0100", B"0111", B"0010", 
 B"0010", B"1001", B"0111", B"1101", 
 B"0101", B"0100", B"0010", B"1000", 
 B"0000", B"1001", B"1011", B"0110", 
 B"1110", B"0100", B"0011", B"1100", 
 B"0001", B"0111", B"0000", B"1001", 
 B"1101", B"0000", B"1111", B"0011", 
 B"1000", B"1011", B"0001", B"0101", 
 B"0001", B"1110", B"1100", B"0101", 
 B"1110", B"0110", B"0011", B"0100", 
 B"0101", B"1111", B"0110", B"0101", 
 B"0011", B"1011", B"0100", B"1110", 
 B"0110", B"1100", B"1010", B"0111", 
 B"1111", B"1100", B"0011", B"1011", 
 B"1101", B"1101", B"1011", B"1011", 
 B"1100", B"0101", B"0001", B"1000", 
 B"1101", B"1100", B"1100", B"0001", 
 B"1101", B"1110", B"0101", B"0110", 
 B"0010", B"1000", B"1100", B"1101", 
 B"0101", B"1001", B"0110", B"1000", 
 B"1011", B"0100", B"0001", B"0100", 
 B"1111", B"1110", B"1000", B"1000", 
 B"0000", B"0001", B"1100", B"1100", 
 B"0101", B"1001", B"1001", B"1101", 
 B"0000", B"0010", B"1001", B"0001", 
 B"1001", B"0111", B"1111", B"1101", 
 B"0001", B"0010", B"0011", B"0010", 
 B"0001", B"0110", B"1111", B"0010", 
 B"0001", B"1000", B"1011", B"1010", 
 B"0100", B"1001", B"0100", B"1110", 
 B"1010", B"1000", B"1100", B"0010", 
 B"1100", B"0101", B"1100", B"1111", 
 B"0100", B"1011", B"0000", B"0101", 
 B"0111", B"0001", B"0110", B"0101", 
 B"0110", B"1011", B"1111", B"1101", 
 B"0111", B"1010", B"0110", B"0011", 
 B"0000", B"0001", B"0101", B"1001", 
 B"1001", B"1001", B"0001", B"1100", 
 B"1010", B"0110", B"0011", B"1111", 
 B"0010", B"1001", B"1110", B"1111", 
 B"0000", B"1011", B"0110", B"1001", 
 B"1101", B"0011", B"0010", B"1100", 
 B"1101", B"1000", B"0001", B"0011", 
 B"0101", B"0110", B"1001", B"0111", 
 B"1010", B"0010", B"1000", B"0100", 
 B"1111", B"0010", B"0000", B"0011", 
 B"1010", B"1010", B"1101", B"0111", 
 B"1011", B"0011", B"0100", B"1111", 
 B"1110", B"0111", B"0111", B"0010", 
 B"0011", B"0111", B"1100", B"0010", 
 B"0101", B"1010", B"0110", B"1111", 
 B"1101", B"0101", B"1100", B"1011", 
 B"1011", B"1011", B"1110", B"0100", 
 B"0111", B"0010", B"1100", B"1101", 
 B"1000", B"0000", B"0110", B"1011", 
 B"0011", B"0001", B"1111", B"0010", 
 B"1101", B"0001", B"0101", B"0111", 
 B"1000", B"1010", B"0000", B"1110", 
 B"1111", B"1111", B"1111", B"1011", 
 B"1110", B"1011", B"1111", B"0001", 
 B"1001", B"0101", B"0011", B"0001", 
 B"0110", B"1001", B"0010", B"0111", 
 B"1111", B"1101", B"1110", B"0110", 
 B"1010", B"1110", B"1100", B"1100", 
 B"1110", B"1111", B"0001", B"1010", 
 B"0111", B"0111", B"1011", B"1000", 
 B"1011", B"0000", B"0011", B"0100", 
 B"1001", B"0110", B"0010", B"1000", 
 B"0001", B"1101", B"1101", B"1010", 
 B"0001", B"1100", B"0000", B"1101", 
 B"0010", B"1111", B"1001", B"1000", 
 B"0100", B"1111", B"0111", B"1011", 
 B"0110", B"0000", B"0001", B"0010", 
 B"1101", B"0110", B"0110", B"0101", 
 B"1111", B"0011", B"1110", B"0101", 
 B"1010", B"1100", B"0101", B"1100", 
 B"0110", B"0010", B"0001", B"0000", 
 B"1101", B"1001", B"0001", B"0100", 
 B"1110", B"1000", B"0110", B"1100", 
 B"1000", B"1100", B"0111", B"1001", 
 B"1001", B"0110", B"1010", B"0001", 
 B"0110", B"0001", B"0101", B"1000", 
 B"0101", B"0101", B"0111", B"0000", 
 B"0111", B"1101", B"0010", B"0001", 
 B"0100", B"0011", B"1110", B"0100", 
 B"1110", B"1000", B"0110", B"1001", 
 B"1101", B"0100", B"0111", B"1000", 
 B"1011", B"0010", B"0111", B"0010", 
 B"1000", B"0110", B"0000", B"1000", 
 B"0101", B"1101", B"0010", B"1100", 
 B"1010", B"0000", B"1111", B"1001", 
 B"0000", B"1001", B"0101", B"0111", 
 B"1000", B"1100", B"0010", B"0001", 
 B"0010", B"1011", B"1000", B"0010", 
 B"0000", B"0100", B"0010", B"0001", 
 B"0100", B"1011", B"0001", B"1100", 
 B"1100", B"0110", B"1001", B"0100", 
 B"0101", B"1110", B"1010", B"0001", 
 B"0110", B"0100", B"1110", B"0111", 
 B"1111", B"1110", B"0001", B"1100", 
 B"0101", B"0000", B"1100", B"0011", 
 B"1001", B"0101", B"0101", B"1100", 
 B"0000", B"0100", B"1011", B"1011", 
 B"0001", B"1011", B"1001", B"1111", 
 B"0100", B"1001", B"0011", B"0000", 
 B"1010", B"1000", B"0110", B"1000", 
 B"0000", B"1101", B"0100", B"1100", 
 B"1110", B"0001", B"0111", B"0001", 
 B"0101", B"0001", B"0101", B"1000", 
 B"1111", B"1000", B"0111", B"1100", 
 B"0111", B"1010", B"0011", B"0010", 
 B"1101", B"0011", B"1011", B"0100", 
 B"1111", B"1101", B"1100", B"1000", 
 B"0100", B"1001", B"0011", B"1110", 
 B"0101", B"0101", B"1100", B"1111", 
 B"1100", B"1100", B"0001", B"1110", 
 B"1000", B"0101", B"1111", B"0101", 
 B"1011", B"1101", B"1001", B"1011", 
 B"1111", B"0001", B"0101", B"0001", 
 B"1000", B"1100", B"0110", B"1010", 
 B"1000", B"0011", B"1111", B"0011", 
 B"1100", B"1101", B"1101", B"1011", 
 B"0000", B"0011", B"1000", B"0001", 
 B"0011", B"1010", B"1000", B"0000", 
 B"0000", B"0111", B"1101", B"1100", 
 B"1110", B"1111", B"0010", B"0100", 
 B"1101", B"1000", B"1010", B"1011", 
 B"1001", B"0010", B"1111", B"1011", 
 B"0111", B"1010", B"1001", B"1110", 
 B"1110", B"0110", B"1101", B"1001", 
 B"0101", B"0101", B"1101", B"1001", 
 B"0101", B"0011", B"1001", B"0101", 
 B"0110", B"1111", B"1101", B"0100", 
 B"1111", B"1011", B"1001", B"1001", 
 B"0111", B"1010", B"0101", B"0010", 
 B"1000", B"1011", B"0100", B"0111", 
 B"0011", B"1101", B"1110", B"0001", 
 B"0101", B"0011", B"1000", B"1101", 
 B"0001", B"0000", B"0111", B"1010", 
 B"1000", B"0010", B"0000", B"0011", 
 B"0100", B"0100", B"0000", B"0111", 
 B"1000", B"0101", B"1001", B"1111", 
 B"1110", B"0010", B"0010", B"0000", 
 B"1100", B"0010", B"0111", B"0000", 
 B"1011", B"1110", B"1101", B"1110", 
 B"0000", B"0010", B"1001", B"0011", 
 B"1111", B"1100", B"0000", B"0101", 
 B"1101", B"0001", B"1110", B"0001", 
 B"1101", B"0000", B"0010", B"0110", 
 B"0000", B"0010", B"0011", B"0100", 
 B"1000", B"1011", B"0001", B"1101", 
 B"1110", B"1000", B"0001", B"0011", 
 B"0100", B"1001", B"0101", B"1001", 
 B"0010", B"1010", B"0001", B"0000", 
 B"1010", B"1110", B"0111", B"1101", 
 B"1111", B"1111", B"0100", B"1111", 
 B"1101", B"1110", B"0101", B"0111", 
 B"0011", B"1101", B"1100", B"1011", 
 B"1110", B"1110", B"0001", B"0101", 
 B"1110", B"1000", B"0111", B"0010", 
 B"0110", B"0111", B"1011", B"0100", 
 B"1110", B"0010", B"0001", B"1110", 
 B"0110", B"1010", B"0101", B"1000", 
 B"0110", B"1010", B"0101", B"1100", 
 B"0001", B"1001", B"1110", B"1000", 
 B"1000", B"1110", B"0101", B"0000", 
 B"1000", B"1101", B"1101", B"0101", 
 B"0001", B"1100", B"1101", B"1110", 
 B"0100", B"1101", B"0100", B"1011", 
 B"0010", B"1110", B"1100", B"0110", 
 B"1101", B"0001", B"0111", B"0001", 
 B"0100", B"0110", B"0100", B"0110", 
 B"1110", B"1011", B"1010", B"0100", 
 B"1011", B"0110", B"1010", B"0010", 
 B"1100", B"1110", B"0011", B"0010", 
 B"1100", B"0110", B"0011", B"1110", 
 B"1010", B"0111", B"0111", B"0010", 
 B"1101", B"1000", B"1111", B"1010", 
 B"1101", B"1001", B"1101", B"0110", 
 B"1010", B"0011", B"0010", B"1001", 
 B"0000", B"0101", B"0100", B"1010", 
 B"1110", B"1001", B"0110", B"1011", 
 B"1000", B"1101", B"1010", B"0010", 
 B"1111", B"1000", B"1011", B"0110", 
 B"1000", B"1010", B"0010", B"1100", 
 B"0000", B"1001", B"0110", B"1111", 
 B"1000", B"0100", B"1111", B"1101", 
 B"1011", B"0000", B"1010", B"0001", 
 B"0011", B"1011", B"1011", B"0010", 
 B"0110", B"1010", B"1000", B"1110", 
 B"0101", B"1010", B"1100", B"1010", 
 B"1110", B"1101", B"0001", B"0101", 
 B"0001", B"0110", B"1101", B"0111", 
 B"1100", B"1111", B"1111", B"0011", 
 B"0111", B"0000", B"0110", B"0100", 
 B"1001", B"1001", B"0100", B"0010", 
 B"1011", B"0010", B"1101", B"0000", 
 B"1110", B"0110", B"1111", B"1101", 
 B"0011", B"0111", B"1100", B"1110", 
 B"1011", B"1101", B"0001", B"1101", 
 B"0011", B"0010", B"1011", B"0011", 
 B"0001", B"1100", B"0001", B"1011", 
 B"0111", B"0101", B"1010", B"1010", 
 B"0001", B"0011", B"1110", B"0000", 
 B"1100", B"0111", B"0001", B"1000", 
 B"0010", B"0000", B"1111", B"0010", 
 B"1110", B"0111", B"1101", B"0011", 
 B"1101", B"1001", B"0001", B"0111", 
 B"1011", B"0101", B"0111", B"0010", 
 B"0100", B"0011", B"1011", B"1110", 
 B"1110", B"1111", B"1101", B"1110", 
 B"1001", B"1011", B"0100", B"0011", 
 B"1001", B"0011", B"1111", B"0100", 
 B"1000", B"1110", B"1001", B"1111", 
 B"1110", B"1100", B"1011", B"0111", 
 B"1001", B"0000", B"0100", B"1010", 
 B"0101", B"0010", B"1001", B"0110", 
 B"0111", B"1111", B"0111", B"0110", 
 B"1000", B"1101", B"0011", B"0111", 
 B"1101", B"1011", B"0000", B"0000", 
 B"1101", B"0100", B"1110", B"0110", 
 B"1010", B"0100", B"1111", B"1010", 
 B"1101", B"1101", B"0110", B"1100"

);

signal data_in          : bit_vector (3 downto 0);
signal reference_data   : bit_vector (3 downto 0);
signal senddata_counter : integer range 0 to 2499 := 2497;

begin

data_in        <= (y0 & y1 & y2 & y3);
senddata       <= senddata_tbl(senddata_counter);
reference_data <= senddata_tbl(senddata_counter);

process (start, clear)
begin
if (clear = '1') then
  senddata_counter <= 2497;
elsif (start = '0' and start'event) then
  if (senddata_counter < 2499) then
     senddata_counter <= senddata_counter + 1;
  else
     senddata_counter <= 0;
  end if;
end if;
end process;

match <= not(data_in xor reference_data);

end verify;
