-- $Id: input.vhdl,v 1.1 2006-01-16 03:40:22 arif_endro Exp $
-------------------------------------------------------------------------------
-- Title       :
-- Project     : 
-------------------------------------------------------------------------------
-- File        :
-- Author      : "Arif E. Nugroho" <arif_endro@yahoo.com>
-- Created     : 2005/12/18
-- Last update : 
-- Simulators  :
-- Synthesizers: ISE Xilinx 6.3i
-- Target      : 
-------------------------------------------------------------------------------
-- Description : 
-------------------------------------------------------------------------------
-- Copyright (C) 2005 Arif E. Nugroho
-- This VHDL design file is an open design; you can redistribute it and/or
-- modify it and/or implement it after contacting the author
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- 
-- 	THIS SOURCE FILE MAY BE USED AND DISTRIBUTED WITHOUT RESTRICTION
-- PROVIDED THAT THIS COPYRIGHT STATEMENT IS NOT REMOVED FROM THE FILE AND THAT
-- ANY DERIVATIVE WORK CONTAINS THE ORIGINAL COPYRIGHT NOTICE AND THE
-- ASSOCIATED DISCLAIMER.
-- 
-------------------------------------------------------------------------------
-- 
-- 	THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY EXPRESS OR
-- IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
-- MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.  IN NO
-- EVENT SHALL THE AUTHOR BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
-- SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
-- PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
-- OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,
-- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR
-- OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity input is
   port (
      clock   : in  bit;
      clear   : in  bit;
      start   : out bit;
      rom_pos : out integer;
      rxin    : out bit_vector (07 downto 00)
      );
end input;

architecture test_bench of input is

type rom_bank is array ( 00000 to 19999 ) of bit_vector (7 downto 0);

constant input_bank : rom_bank :=
(

 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"00100000", B"00100000", B"11100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"00100000", B"00100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"00100000",
 B"00100000", B"11100000", B"11100000", B"11100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"00100000", B"00100000",
 B"11100000", B"00100000", B"11100000", B"00100000", B"11100000",
 B"11100000", B"00100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"11100000",
 B"00100000", B"11100000", B"11100000", B"00100000", B"00100000",
 B"11100000", B"11100000", B"00100000", B"11100000", B"11100000",
 B"11100000", B"11100000", B"11100000", B"11100000", B"00100000",
 B"00100000", B"00100000", B"00100000", B"11100000", B"11100000"

);

signal input_counter : integer range 0 to 19999 := 0;
signal start_fifo    : bit_vector (7 downto 0) := ( B"0100_0000" );
signal clk : bit;

begin

process (clk, clear)
begin
if (clear = '1') then
    rxin <= (others => '0');
elsif (clk = '1' and clk'event) then
    rxin <= input_bank(input_counter);
end if;
end process;

process (clk, clear)
begin
if (clear = '1') then
    input_counter <= 0;
elsif (clk = '1' and clk'event) then
    if (input_counter < 19999) then
    input_counter <= input_counter + 1;
    else
    input_counter <= 0;
    end if;
end if;
end process;

rom_pos <= input_counter;

process (clk, clear)
begin
if (clear = '1') then
    start_fifo <= B"0100_0000";
elsif ( clk = '1' and clk'event) then
    start_fifo <= start_fifo (6 downto 0) & start_fifo (7);
end if;
end process;

clk   <= clock;
start <= start_fifo (7);

end test_bench;
