-- $Id: input6DB.vhdl,v 1.1 2006-01-16 03:40:22 arif_endro Exp $
-------------------------------------------------------------------------------
-- Title       :
-- Project     : 
-------------------------------------------------------------------------------
-- File        :
-- Author      : "Arif E. Nugroho" <arif_endro@yahoo.com>
-- Created     : 2005/12/18
-- Last update : 
-- Simulators  :
-- Synthesizers: ISE Xilinx 6.3i
-- Target      : 
-------------------------------------------------------------------------------
-- Description : 
-------------------------------------------------------------------------------
-- Copyright (C) 2005 Arif E. Nugroho
-- This VHDL design file is an open design; you can redistribute it and/or
-- modify it and/or implement it after contacting the author
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- 
-- 	THIS SOURCE FILE MAY BE USED AND DISTRIBUTED WITHOUT RESTRICTION
-- PROVIDED THAT THIS COPYRIGHT STATEMENT IS NOT REMOVED FROM THE FILE AND THAT
-- ANY DERIVATIVE WORK CONTAINS THE ORIGINAL COPYRIGHT NOTICE AND THE
-- ASSOCIATED DISCLAIMER.
-- 
-------------------------------------------------------------------------------
-- 
-- 	THIS SOFTWARE IS PROVIDED BY THE AUTHOR ``AS IS'' AND ANY EXPRESS OR
-- IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF
-- MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.  IN NO
-- EVENT SHALL THE AUTHOR BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
-- SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
-- PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
-- OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY,
-- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR
-- OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity input is
   port (
      clock   : in  bit;
      clear   : in  bit;
      start   : out bit;
      rom_pos : out integer;
      rxin    : out bit_vector (07 downto 00)
      );
end input;

architecture test_bench of input is

type rom_bank is array ( 00000 to 19999 ) of bit_vector (7 downto 0);

constant input_bank : rom_bank :=
(

 B"00110111", B"00100110", B"11100011", B"00101110", B"00100101",
 B"11100111", B"11110011", B"00011110", B"00101100", B"00100001",
 B"00010111", B"11010110", B"00110010", B"11100101", B"00000001",
 B"11010110", B"11011110", B"11011101", B"00010100", B"11010011",
 B"00001001", B"11011110", B"10101000", B"00010011", B"11010110",
 B"00011111", B"11011011", B"11101001", B"11101100", B"00110111",
 B"00100101", B"11010110", B"11101101", B"00010111", B"00011001",
 B"00010010", B"11100110", B"00100010", B"11101001", B"00101101",
 B"11111000", B"00101000", B"11010110", B"11100110", B"11010110",
 B"00010001", B"00011001", B"00001001", B"11000110", B"11110000",
 B"00011110", B"11001101", B"00100011", B"11001011", B"11100101",
 B"00001011", B"11010100", B"11111001", B"00101110", B"00001011",
 B"00101000", B"00010010", B"11101000", B"11100000", B"00100101",
 B"00011010", B"11100100", B"00010010", B"00100101", B"11100001",
 B"11010111", B"00100110", B"00100001", B"00010101", B"11101011",
 B"11101110", B"00111011", B"00000110", B"11110010", B"11101100",
 B"11011111", B"00000101", B"00001110", B"00000100", B"00100110",
 B"00011010", B"11110011", B"11111001", B"11000111", B"00111010",
 B"11101000", B"00011010", B"11100101", B"11101101", B"00011011",
 B"00001101", B"11101101", B"00001011", B"00110000", B"11101111",
 B"11001110", B"11011100", B"11011000", B"11000110", B"11100111",
 B"11010010", B"11001100", B"11011110", B"00011100", B"00010110",
 B"00001110", B"00010000", B"00011111", B"11100011", B"11001010",
 B"00010110", B"11100111", B"11010100", B"11101010", B"11111111",
 B"00000010", B"00110000", B"11100101", B"00010100", B"00100101",
 B"11101000", B"11010010", B"00011100", B"11100101", B"11100000",
 B"00101100", B"00011000", B"00110010", B"00001010", B"11011101",
 B"11010111", B"11101100", B"00100111", B"00010110", B"00010011",
 B"11111001", B"00011000", B"11111000", B"00001000", B"00010101",
 B"00001110", B"00100011", B"11101111", B"00010010", B"11011001",
 B"00101101", B"11001101", B"11011111", B"00011010", B"11001011",
 B"01001011", B"11011100", B"11011000", B"00100000", B"00100011",
 B"00010111", B"11011110", B"11100111", B"00011001", B"11010110",
 B"11001011", B"11110110", B"11110100", B"11010110", B"00001101",
 B"11011100", B"00000001", B"11101111", B"00001010", B"00001010",
 B"11011110", B"01000010", B"11010101", B"00110100", B"11010011",
 B"11101111", B"11001100", B"00011110", B"00010001", B"00101001",
 B"00010100", B"00101111", B"11011000", B"00010111", B"11100011",
 B"00110010", B"11110010", B"11101111", B"11100110", B"00111001",
 B"00110111", B"00100110", B"00010100", B"11100010", B"11100010",
 B"11001010", B"00100100", B"00101000", B"11011000", B"11011010",
 B"11011100", B"11110000", B"11101000", B"11010101", B"11110111",
 B"00001000", B"00001101", B"00010110", B"01001011", B"11011001",
 B"11111011", B"11011000", B"00011110", B"00010101", B"00100010",
 B"11010110", B"00010110", B"11000100", B"00001101", B"00110010",
 B"11010110", B"11010110", B"00011001", B"11100100", B"11011100",
 B"11100011", B"11011001", B"11101110", B"11101101", B"00011000",
 B"11011101", B"00110010", B"11011101", B"11011100", B"00010111",
 B"00010011", B"00100011", B"00100110", B"00110111", B"00011101",
 B"00011011", B"00100010", B"00010001", B"00010100", B"11011001",
 B"00011101", B"00110100", B"11010101", B"00110010", B"00110001",
 B"11011101", B"00100111", B"00000010", B"00001001", B"00100101",
 B"00011001", B"00100010", B"00100010", B"00000001", B"00010111",
 B"11000110", B"11010110", B"00010001", B"11101000", B"11010110",
 B"11101110", B"11011001", B"11001110", B"11100110", B"00010100",
 B"11111001", B"00010010", B"11110111", B"11100010", B"00001101",
 B"11111001", B"00011001", B"11111110", B"11100100", B"11010100",
 B"00101011", B"00111101", B"11101101", B"00011001", B"00011000",
 B"00100000", B"00010000", B"00010001", B"00011101", B"00001100",
 B"00001011", B"11000101", B"00011011", B"00110000", B"11011110",
 B"11010000", B"11110001", B"11100101", B"11010111", B"11010001",
 B"00010011", B"00101100", B"11100100", B"11100000", B"11010100",
 B"11100000", B"11111001", B"11011011", B"00101100", B"00011001",
 B"00110011", B"11100110", B"00010001", B"11010011", B"00011011",
 B"00101001", B"11101001", B"11010001", B"00100111", B"11011011",
 B"11111101", B"11100100", B"11110001", B"11110111", B"11011101",
 B"00100100", B"00010101", B"00100111", B"00001010", B"11011011",
 B"11010111", B"00011111", B"11010101", B"11101001", B"00100100",
 B"11110110", B"11110000", B"11001011", B"11010011", B"11110000",
 B"11010010", B"00011111", B"11111010", B"00011101", B"11100101",
 B"11110001", B"00100110", B"11110111", B"11101001", B"00001000",
 B"11010111", B"00001001", B"11110010", B"11010001", B"00010111",
 B"11010101", B"00001100", B"11100111", B"11001110", B"11010100",
 B"00101000", B"00011001", B"11110000", B"00010000", B"11011101",
 B"00100010", B"11011110", B"11011011", B"11101010", B"00110000",
 B"00011101", B"11100001", B"11011110", B"00100100", B"11010000",
 B"00100011", B"11011010", B"11101110", B"00101011", B"11100011",
 B"11011111", B"11010101", B"11011010", B"00010110", B"00101011",
 B"00101010", B"00011101", B"00011000", B"11110011", B"11101000",
 B"00111111", B"11110010", B"11100010", B"11100000", B"11110111",
 B"11100101", B"00010100", B"00011011", B"00100110", B"11010010",
 B"00110010", B"11101010", B"00011101", B"00110001", B"00110001",
 B"11010101", B"00101001", B"00100111", B"11101111", B"11001001",
 B"11110100", B"00000010", B"11011000", B"11111100", B"11110110",
 B"00101010", B"00010101", B"00100110", B"00110000", B"00110101",
 B"11100010", B"11001001", B"00101101", B"11101111", B"11100111",
 B"11000011", B"11001101", B"00011100", B"00010110", B"00100000",
 B"00010000", B"00101011", B"00100000", B"00111001", B"00100110",
 B"11101111", B"11101110", B"11011011", B"00011100", B"00100111",
 B"11110111", B"00100010", B"11010001", B"00010010", B"00110000",
 B"00110100", B"11111000", B"00011000", B"11101111", B"00100000",
 B"11111001", B"00101111", B"11010001", B"00111001", B"11001100",
 B"11010010", B"11011100", B"00011000", B"00101010", B"00110110",
 B"11010100", B"11010010", B"11011001", B"11001111", B"00100011",
 B"11111000", B"00110011", B"11011010", B"10111100", B"11011111",
 B"11011110", B"00011110", B"00011111", B"00011010", B"00101100",
 B"00100010", B"00000010", B"00010101", B"00011000", B"11101100",
 B"00100111", B"00011110", B"11010011", B"11000111", B"00010000",
 B"11011001", B"00101001", B"11010101", B"11000010", B"00011110",
 B"00110010", B"11101100", B"00111010", B"11101011", B"11010100",
 B"10111101", B"00001010", B"00010010", B"11011100", B"00101111",
 B"11101101", B"11010000", B"11101011", B"11011010", B"00111110",
 B"11100001", B"00110000", B"00011000", B"00101100", B"11011000",
 B"11100000", B"00100011", B"00101110", B"11000110", B"11100110",
 B"11100100", B"11110100", B"00100010", B"11100000", B"00101100",
 B"11011110", B"11001000", B"00100010", B"11010110", B"00101111",
 B"00111010", B"00110001", B"11010110", B"00100000", B"11010010",
 B"00010100", B"11101100", B"00010101", B"00100101", B"00100111",
 B"11100110", B"00100100", B"11110011", B"00011111", B"00111001",
 B"00001101", B"00010100", B"10111111", B"00011010", B"11110011",
 B"00001111", B"11010010", B"11101001", B"01000001", B"00111111",
 B"11111101", B"11100110", B"00110100", B"11001111", B"00011010",
 B"11100110", B"11001001", B"11001100", B"00101000", B"01000010",
 B"11001000", B"00101001", B"11010010", B"00011100", B"11010111",
 B"11100001", B"00111000", B"11001000", B"11100101", B"11000101",
 B"11010011", B"11010010", B"11010010", B"11010010", B"11100001",
 B"01000011", B"00001001", B"00101101", B"00010011", B"11110011",
 B"11010100", B"00101001", B"11011011", B"00011000", B"11111000",
 B"11010010", B"00011110", B"00110101", B"00001111", B"00100101",
 B"00011101", B"00100011", B"11111111", B"00011010", B"00100001",
 B"00110111", B"00110100", B"00011011", B"00001001", B"00100100",
 B"00101101", B"00101011", B"00100101", B"11100110", B"11010110",
 B"00000100", B"11010000", B"00101100", B"00100001", B"00101101",
 B"00110000", B"11100110", B"00010111", B"11100000", B"11101101",
 B"11010010", B"11101001", B"00101010", B"00100111", B"11011000",
 B"00010011", B"00011011", B"11000111", B"11010100", B"11011101",
 B"11101011", B"11000001", B"01000111", B"00100101", B"00001011",
 B"11100110", B"00100110", B"00100111", B"11011110", B"00010000",
 B"11110100", B"11011100", B"11100111", B"00100101", B"00100010",
 B"00000111", B"00000101", B"11101001", B"00101111", B"00011101",
 B"11101100", B"00001101", B"00100100", B"11011000", B"11100110",
 B"00110111", B"00001110", B"00001011", B"11000111", B"00001010",
 B"00010110", B"11001000", B"11011011", B"00101101", B"00100101",
 B"00010111", B"11010101", B"11101111", B"00100000", B"00101000",
 B"11011010", B"11011110", B"00000101", B"00010010", B"00100011",
 B"00010101", B"11001000", B"00100010", B"11110011", B"00011001",
 B"11011100", B"11100000", B"00101010", B"11100010", B"00100001",
 B"11000111", B"11101010", B"00110011", B"11100001", B"11000101",
 B"00010110", B"11111100", B"00010110", B"11100110", B"11101000",
 B"00101111", B"00100100", B"00101011", B"00010100", B"00100010",
 B"00101011", B"00110100", B"00011100", B"00110110", B"00011011",
 B"00001110", B"00011010", B"00001011", B"00100001", B"00010100",
 B"00101100", B"00011011", B"11010011", B"00101001", B"00010101",
 B"11100111", B"11101001", B"11100111", B"11110101", B"11101111",
 B"11001001", B"00100110", B"11010100", B"00001010", B"11101000",
 B"00001111", B"00100000", B"00101011", B"11110100", B"00100011",
 B"11100100", B"00101101", B"11110010", B"11011100", B"00100010",
 B"00101000", B"00100111", B"00100100", B"00110010", B"00100011",
 B"00010111", B"00110000", B"00011001", B"00100110", B"00101000",
 B"11101110", B"11001111", B"11100010", B"11011001", B"00100111",
 B"11010000", B"00101011", B"00011001", B"00110001", B"00011000",
 B"11001101", B"00100100", B"11011111", B"00010111", B"11011111",
 B"11010111", B"11011111", B"11011010", B"11101010", B"00110000",
 B"00101110", B"00101101", B"00010000", B"11100100", B"00001000",
 B"11000111", B"00110001", B"11000101", B"11010011", B"01000110",
 B"00101110", B"00110101", B"10110100", B"11100100", B"00000111",
 B"11110000", B"11100001", B"11100101", B"11011100", B"00011101",
 B"11101000", B"00000001", B"00111001", B"11111111", B"11111100",
 B"00100101", B"11111111", B"00100010", B"00001001", B"00011001",
 B"00101000", B"00011000", B"00011010", B"11111110", B"00001110",
 B"11101101", B"00010110", B"11011101", B"11110000", B"11001000",
 B"00100100", B"00011000", B"11001010", B"11101011", B"11110000",
 B"00011100", B"00111110", B"00110000", B"00001001", B"11010010",
 B"11001100", B"00011010", B"00101010", B"00010011", B"00011111",
 B"00111000", B"00011011", B"00011011", B"00101011", B"00010001",
 B"00010101", B"11010010", B"11010011", B"00110100", B"00001101",
 B"11100001", B"11101011", B"11110010", B"11100100", B"10110110",
 B"11100100", B"00011010", B"00010011", B"00011011", B"00100100",
 B"00000100", B"00111100", B"00010001", B"11100100", B"00001001",
 B"11100001", B"00011110", B"11100000", B"00101100", B"00101001",
 B"00001111", B"00101000", B"00001001", B"00011001", B"00010000",
 B"00010111", B"00011111", B"00011011", B"00101101", B"00010110",
 B"00001010", B"00001100", B"00101010", B"00100011", B"11100011",
 B"00001111", B"11111110", B"10111110", B"11110010", B"00101111",
 B"00101001", B"11111110", B"00100000", B"11110010", B"00100001",
 B"00100100", B"11110000", B"00011010", B"00100101", B"11011110",
 B"11011011", B"11101101", B"00100000", B"11001000", B"00010111",
 B"11101110", B"11011001", B"11110111", B"00110011", B"00010001",
 B"11010100", B"10110011", B"00100010", B"11111110", B"11101011",
 B"11010001", B"11111101", B"00001000", B"00101001", B"11010010",
 B"00110110", B"11010101", B"00000101", B"11001101", B"11010110",
 B"00101101", B"01000001", B"00101110", B"11101011", B"00100111",
 B"11001001", B"00100001", B"00011101", B"11010011", B"00110001",
 B"11100100", B"11101001", B"11101111", B"00010101", B"00100110",
 B"00011011", B"00100000", B"00100011", B"00101111", B"00100001",
 B"00011110", B"00110111", B"00010000", B"00111011", B"11110101",
 B"00011010", B"00100111", B"11010101", B"00011110", B"00000101",
 B"11000111", B"11011101", B"11001101", B"11010100", B"11011111",
 B"00011101", B"00011100", B"00101010", B"00101010", B"00100111",
 B"11101110", B"00010110", B"00100101", B"11100100", B"00011111",
 B"00101110", B"11100110", B"00100100", B"00101111", B"11101101",
 B"00110100", B"00100101", B"11100110", B"11011000", B"00011010",
 B"00101100", B"11110010", B"00101100", B"11010001", B"11110000",
 B"11011100", B"00100011", B"00001100", B"00100001", B"00010111",
 B"01000010", B"00100010", B"00100000", B"00011001", B"11110011",
 B"00100011", B"00101010", B"00011010", B"00101001", B"11110111",
 B"00100000", B"11101000", B"00011001", B"11110101", B"01000111",
 B"11100001", B"00100001", B"00110010", B"11011000", B"00001011",
 B"00010110", B"11100011", B"11011001", B"00010110", B"00000101",
 B"00101000", B"11100110", B"00100001", B"11110010", B"00011110",
 B"01001011", B"00000110", B"00000000", B"00001000", B"00011111",
 B"00100010", B"00011000", B"00100000", B"11111001", B"11100000",
 B"00101111", B"11011111", B"00010010", B"11100100", B"11010000",
 B"00010111", B"11101000", B"11100110", B"00110011", B"00100111",
 B"00101011", B"00100101", B"11010010", B"11100101", B"10111001",
 B"11011100", B"00000011", B"00101111", B"00101001", B"11110001",
 B"00010011", B"11101010", B"11101110", B"11110100", B"00110000",
 B"00011100", B"00000000", B"00100101", B"11100001", B"11110111",
 B"11011101", B"00100000", B"00101100", B"11100010", B"11011101",
 B"11100001", B"11111011", B"11010111", B"00011100", B"00010011",
 B"11100001", B"00100001", B"00001010", B"11010000", B"11111111",
 B"00100110", B"00001101", B"11110001", B"11111110", B"11101111",
 B"11100101", B"11011001", B"00100001", B"00100010", B"00101100",
 B"00011010", B"00011001", B"11011010", B"00001101", B"11101001",
 B"00011100", B"11101001", B"00100011", B"11110011", B"00001101",
 B"11011011", B"11100111", B"11010011", B"00010101", B"00011100",
 B"11001011", B"00001100", B"00010111", B"11001100", B"11101110",
 B"11010111", B"11101101", B"10111110", B"00100000", B"00101111",
 B"11011000", B"11100001", B"00100100", B"00000110", B"11101001",
 B"11010000", B"11011000", B"00011101", B"11011010", B"00110011",
 B"11100001", B"11110100", B"00011000", B"00001111", B"00011101",
 B"11010010", B"11101000", B"11001110", B"11001111", B"00101011",
 B"11100000", B"00001001", B"11110010", B"11100110", B"00011010",
 B"11101111", B"00110110", B"10110100", B"10111101", B"00100010",
 B"00101101", B"00010110", B"10110011", B"00010010", B"00101000",
 B"11001011", B"11110000", B"00010111", B"11001011", B"11110000",
 B"11011111", B"11010101", B"11111110", B"01000100", B"00010110",
 B"00100100", B"11010011", B"00100000", B"11101101", B"00010000",
 B"11001011", B"11100011", B"00011000", B"00010001", B"00010010",
 B"00011011", B"11110001", B"11101000", B"01000110", B"00010011",
 B"11000100", B"11100001", B"00100000", B"00011011", B"11100001",
 B"11100001", B"00110100", B"00010110", B"11011111", B"11001100",
 B"00100000", B"00100001", B"11010100", B"00000110", B"00100010",
 B"11110010", B"11100111", B"00001100", B"00100100", B"11001100",
 B"11100111", B"11111011", B"11001100", B"00101000", B"11110110",
 B"00010001", B"00011011", B"00000100", B"11101111", B"00110000",
 B"00001011", B"11100010", B"11100011", B"00101100", B"00011010",
 B"00011100", B"00000101", B"00010010", B"00010111", B"00100001",
 B"00110000", B"00010100", B"00101001", B"00101011", B"00001010",
 B"11011111", B"00100000", B"11110011", B"00100010", B"11001001",
 B"00000001", B"11101111", B"11100111", B"00001110", B"11100011",
 B"11011001", B"11011111", B"11011010", B"11100100", B"11011001",
 B"00101110", B"00011100", B"00101010", B"00001000", B"11101100",
 B"00001010", B"00000110", B"00010000", B"00010011", B"11010100",
 B"00100100", B"11101000", B"00100110", B"11011100", B"00011101",
 B"00000110", B"11101010", B"00100100", B"11100000", B"11101111",
 B"11010001", B"11000101", B"11100011", B"11110001", B"11110101",
 B"00011101", B"00101000", B"11100100", B"00001100", B"11000111",
 B"00011010", B"11011110", B"11100101", B"11111100", B"11010010",
 B"11111000", B"11101101", B"11000101", B"11100010", B"11001011",
 B"00101011", B"11100011", B"00101010", B"11101011", B"11011000",
 B"00001111", B"00101010", B"00011100", B"00000110", B"11011011",
 B"00011101", B"11101101", B"00000001", B"11001111", B"11101001",
 B"11011001", B"00100110", B"00000000", B"00011010", B"11010111",
 B"11001010", B"00101010", B"00101001", B"00100001", B"00101111",
 B"11011011", B"00001001", B"11010100", B"00011101", B"11110000",
 B"00110010", B"01000001", B"00001101", B"11101011", B"01001011",
 B"00110110", B"10110000", B"11101100", B"11011111", B"00101000",
 B"00110000", B"00010001", B"11001100", B"00111110", B"11010111",
 B"00000101", B"11011100", B"00011001", B"00001111", B"11011111",
 B"11011111", B"11010010", B"11000010", B"11001010", B"11100100",
 B"00110001", B"11001100", B"00010001", B"11101100", B"11011110",
 B"00101110", B"00010000", B"00100010", B"11011100", B"11100010",
 B"01000011", B"11101011", B"11011000", B"11010111", B"11001101",
 B"11101110", B"11010110", B"00001011", B"11101010", B"00111111",
 B"11101000", B"11001101", B"00000001", B"00110001", B"11011010",
 B"11010110", B"00000111", B"11010011", B"11011011", B"11110101",
 B"11110000", B"11011100", B"00010000", B"11000110", B"00110010",
 B"11011100", B"11001011", B"11110111", B"00011011", B"00110011",
 B"00100101", B"00000000", B"11011111", B"01000100", B"00100110",
 B"11011000", B"11011111", B"00010101", B"00011111", B"11111101",
 B"00011110", B"00010100", B"11101100", B"11011110", B"00011001",
 B"11111101", B"11101011", B"11111000", B"00100011", B"00101010",
 B"11011100", B"00010110", B"11101001", B"11010111", B"11110101",
 B"00110000", B"11001010", B"00010000", B"11110010", B"11110100",
 B"00101001", B"11101110", B"00011101", B"11101011", B"11011010",
 B"11011110", B"00010110", B"00100001", B"11011110", B"00111110",
 B"00110010", B"11100010", B"00100001", B"01000100", B"11100010",
 B"11100111", B"00110000", B"11100110", B"11101100", B"11100010",
 B"00110010", B"00100010", B"11100001", B"00110000", B"11100001",
 B"11101000", B"11110010", B"00110011", B"00100101", B"11010011",
 B"00010011", B"11011100", B"00100001", B"00011100", B"00100011",
 B"11011111", B"00010010", B"01001100", B"11100011", B"11100010",
 B"00101010", B"11011110", B"11100010", B"11111000", B"11101100",
 B"00111000", B"00101111", B"00011001", B"11111111", B"00110101",
 B"00010110", B"11011100", B"00101001", B"00011110", B"11011010",
 B"11011000", B"00011111", B"00100001", B"11010001", B"11000111",
 B"00110010", B"11000011", B"11110100", B"11011011", B"11100011",
 B"11010011", B"11011111", B"00000011", B"00101101", B"11111100",
 B"11100011", B"00110000", B"11100101", B"11100110", B"11100001",
 B"00010001", B"00010110", B"01000110", B"00010101", B"11100110",
 B"10110101", B"00101110", B"00010111", B"00100110", B"00001001",
 B"00001010", B"00001111", B"11111110", B"00001100", B"00101110",
 B"00001010", B"11111001", B"00101111", B"00010110", B"00101000",
 B"00010110", B"11111111", B"11111011", B"00010111", B"00011111",
 B"00110110", B"00010110", B"00011011", B"00100111", B"00101111",
 B"00110100", B"11101101", B"11010011", B"00001100", B"10110110",
 B"11001100", B"11101101", B"11101010", B"11110110", B"11101111",
 B"11001100", B"00000101", B"00010101", B"11101011", B"00011001",
 B"11101010", B"00100001", B"11011011", B"00101111", B"11010110",
 B"11100011", B"11100010", B"00001101", B"00111001", B"11110001",
 B"00011000", B"11011101", B"00010010", B"11100100", B"11110101",
 B"00011000", B"00101001", B"11110101", B"00011001", B"00011000",
 B"00101100", B"11010111", B"00100101", B"11000010", B"00011011",
 B"00010110", B"11011100", B"00110011", B"00010010", B"11101001",
 B"00110110", B"00010010", B"11101100", B"00111110", B"00010011",
 B"00010000", B"11110110", B"00010011", B"11100111", B"00110010",
 B"11000101", B"00100100", B"00001000", B"00101000", B"11011010",
 B"11100001", B"11100000", B"00100110", B"00011001", B"00001100",
 B"11010011", B"11010100", B"00010101", B"11100111", B"11111110",
 B"11101100", B"11011111", B"11011100", B"11010110", B"00101101",
 B"11110110", B"00001111", B"11001110", B"11000000", B"00100110",
 B"11110100", B"00100111", B"11100100", B"11011001", B"11101111",
 B"00011111", B"00100100", B"11100110", B"11011011", B"00100010",
 B"00110001", B"00100011", B"11011101", B"00110111", B"11001101",
 B"00101100", B"11101000", B"11100110", B"11011011", B"11110011",
 B"00100000", B"00010101", B"00100110", B"00101011", B"11011111",
 B"11101000", B"11010001", B"11111011", B"00100111", B"00101000",
 B"00101001", B"01000101", B"11110010", B"11010001", B"00011110",
 B"11001111", B"00010000", B"11010100", B"11100111", B"00001100",
 B"00101000", B"00001110", B"00011010", B"11101100", B"00100101",
 B"11011100", B"00100001", B"11100011", B"11011101", B"00101010",
 B"11001110", B"11101001", B"11011011", B"00001110", B"00000111",
 B"11100010", B"11011101", B"00111001", B"00011000", B"00010110",
 B"11010111", B"00101011", B"11000100", B"00110111", B"00111010",
 B"00100011", B"11010011", B"11001100", B"01010100", B"00100111",
 B"11010101", B"11110101", B"00101101", B"00000010", B"11100110",
 B"00111111", B"00011111", B"11111011", B"11011011", B"00100111",
 B"00110000", B"11101101", B"00011000", B"00010011", B"11011000",
 B"00100111", B"00010100", B"11100101", B"00011000", B"00101010",
 B"11001010", B"00001011", B"00100100", B"11000000", B"11001101",
 B"00100010", B"00101001", B"00101110", B"00000100", B"00111111",
 B"00100110", B"11101100", B"11010101", B"00011110", B"00101001",
 B"01001101", B"11110000", B"00111001", B"00100001", B"11110000",
 B"11001111", B"00011010", B"00100000", B"11110011", B"00111010",
 B"11001111", B"11001101", B"11011000", B"00011100", B"00110011",
 B"00011100", B"11011001", B"11011100", B"10111110", B"11110110",
 B"00010011", B"11110011", B"00110011", B"11100000", B"11100111",
 B"00001010", B"11101100", B"00001100", B"11011011", B"11101000",
 B"00010111", B"11011111", B"11111011", B"00001001", B"00110011",
 B"11111001", B"00010110", B"11101001", B"00000110", B"11000110",
 B"11000110", B"00101011", B"11001100", B"00101011", B"11001101",
 B"11001101", B"00010010", B"11011110", B"00010100", B"00011111",
 B"11001101", B"11101111", B"11101011", B"11010101", B"11001001",
 B"11011100", B"00001111", B"00101101", B"11100000", B"11111011",
 B"11001010", B"11110100", B"11101101", B"00011010", B"11001100",
 B"00100111", B"11011000", B"11101101", B"11100110", B"00100001",
 B"00010011", B"00011010", B"00010100", B"11110010", B"11010001",
 B"00010000", B"00011010", B"11110011", B"11101101", B"00101001",
 B"11101111", B"00000110", B"00001111", B"11100101", B"00101001",
 B"00100010", B"11011101", B"00011100", B"00011110", B"00010011",
 B"00010101", B"00011111", B"00101101", B"00011000", B"00100011",
 B"11000110", B"11010101", B"00011110", B"00010111", B"00100001",
 B"00010101", B"11011000", B"11011100", B"11011111", B"11110010",
 B"00101001", B"00100001", B"00101101", B"00100100", B"11010110",
 B"11101011", B"11001010", B"11111101", B"00010111", B"00011001",
 B"11011111", B"00100101", B"11011111", B"00100000", B"11011101",
 B"00101000", B"00100000", B"11101010", B"11100011", B"11100001",
 B"11101111", B"11011111", B"00011110", B"00001011", B"00001111",
 B"00001000", B"00101001", B"00010100", B"00001000", B"00110001",
 B"11100110", B"11011111", B"11110110", B"00001010", B"00101111",
 B"11011010", B"00000010", B"11101001", B"00001001", B"11100101",
 B"11010101", B"00001000", B"11101101", B"11010111", B"11100010",
 B"11100101", B"11011110", B"11011101", B"00010110", B"11001010",
 B"00011001", B"11110101", B"11011110", B"00111011", B"00101100",
 B"00100001", B"11101001", B"00011011", B"00011111", B"11011100",
 B"11011000", B"00100111", B"00011100", B"00111110", B"01000001",
 B"00011100", B"00011101", B"00010011", B"00111110", B"00100110",
 B"11110010", B"11101110", B"11101000", B"10110111", B"00101101",
 B"00110010", B"00110010", B"00101101", B"11001001", B"00000110",
 B"11100101", B"00110101", B"11011010", B"10111101", B"00011011",
 B"00100010", B"11010011", B"00110010", B"11101010", B"00101000",
 B"11011110", B"11101100", B"11111110", B"00111010", B"00111011",
 B"11101001", B"11111010", B"00100110", B"11001010", B"01000001",
 B"00101010", B"11100001", B"11100010", B"11001011", B"00100000",
 B"11011010", B"00010101", B"11100010", B"11100011", B"00101110",
 B"00001111", B"00011111", B"11101110", B"00101101", B"00100010",
 B"11110010", B"11001110", B"00100110", B"11110000", B"00000000",
 B"00110111", B"11010111", B"11110010", B"11011110", B"11100110",
 B"11011000", B"11000100", B"00110110", B"00001001", B"11011011",
 B"11110110", B"11101011", B"11001110", B"11101111", B"11100100",
 B"00001101", B"11011100", B"11100100", B"11011111", B"00101011",
 B"00101000", B"11100001", B"11011001", B"00011001", B"00110011",
 B"00010010", B"11101110", B"00010001", B"11000101", B"11111101",
 B"00001100", B"00001111", B"00101011", B"00010111", B"00011011",
 B"11110111", B"00110010", B"00011010", B"11100010", B"00100111",
 B"00011110", B"11111000", B"11010111", B"11001111", B"11110100",
 B"11010110", B"11000110", B"11100100", B"11110001", B"00101100",
 B"00001010", B"11111110", B"00100100", B"11101100", B"00010011",
 B"00110100", B"00110001", B"00101010", B"00100010", B"00001001",
 B"00100001", B"00001110", B"00100111", B"11111010", B"11010011",
 B"00100010", B"11001110", B"11011000", B"11011110", B"11101110",
 B"11111001", B"00100001", B"00001001", B"00011110", B"11100100",
 B"00100010", B"00010000", B"00110111", B"00101010", B"11011001",
 B"00001111", B"11000011", B"11110101", B"11001101", B"00101001",
 B"00000111", B"11110110", B"00100000", B"11011000", B"00010100",
 B"01000110", B"11001011", B"11011001", B"00001110", B"11011011",
 B"11100010", B"00101001", B"00100011", B"00100010", B"00101000",
 B"11011010", B"11101101", B"01000110", B"11011100", B"00100101",
 B"00010110", B"11001000", B"00100010", B"00101110", B"11001111",
 B"11100110", B"00101010", B"00001100", B"00110101", B"11101101",
 B"00001011", B"11010110", B"00011001", B"00011111", B"11011000",
 B"11001000", B"00010110", B"11100100", B"11011110", B"11111011",
 B"11100101", B"00011000", B"11011100", B"00011001", B"00011111",
 B"11101100", B"00111000", B"00011100", B"11011011", B"11010100",
 B"11100001", B"11110101", B"11110001", B"00100101", B"00011010",
 B"00011000", B"00100100", B"11111000", B"00100010", B"11001000",
 B"11011001", B"00110001", B"00100111", B"11010010", B"11100010",
 B"00100111", B"11101111", B"00010010", B"11101100", B"11100001",
 B"11001010", B"00000001", B"00011101", B"00011010", B"00100010",
 B"00110100", B"00010110", B"00011000", B"00100000", B"00110110",
 B"00101001", B"11010110", B"11011100", B"00011101", B"01000100",
 B"00101100", B"00011110", B"11010101", B"11011100", B"00110011",
 B"11001010", B"11101011", B"00100011", B"11111101", B"11011110",
 B"11010100", B"11111000", B"11011111", B"11101110", B"11010110",
 B"00010110", B"00011100", B"11010111", B"00010011", B"11101010",
 B"11101001", B"11100011", B"11010101", B"11100001", B"00010000",
 B"00100100", B"00100111", B"00010111", B"11000101", B"00111100",
 B"00011101", B"00011010", B"00000000", B"00100011", B"11101101",
 B"00011010", B"11100011", B"00010011", B"00100010", B"00011100",
 B"11011011", B"00010001", B"11001010", B"00010010", B"00010110",
 B"11100000", B"11010111", B"00010000", B"11011001", B"11011101",
 B"11011111", B"11011100", B"11010101", B"00100101", B"00011011",
 B"00011011", B"11101111", B"00011101", B"11100101", B"00101000",
 B"11100011", B"00010101", B"00000100", B"00101110", B"11010111",
 B"00001100", B"11100011", B"00111110", B"11100000", B"11011010",
 B"00110001", B"00101001", B"00011011", B"00100001", B"11010111",
 B"11111101", B"11100001", B"00100001", B"00001000", B"00011100",
 B"11100101", B"00011010", B"11000001", B"00010101", B"11000100",
 B"11110100", B"00100111", B"00001110", B"00100001", B"00000101",
 B"00000011", B"11100011", B"00110100", B"00011100", B"11110000",
 B"11100010", B"00011101", B"00101101", B"11010101", B"11011111",
 B"00011000", B"11001101", B"11100111", B"00011111", B"11101100",
 B"11100111", B"11011011", B"11101110", B"11010100", B"00001000",
 B"00011100", B"11110011", B"11010100", B"11100111", B"11101100",
 B"11010100", B"00101110", B"11101100", B"00011100", B"11100010",
 B"11010110", B"11110001", B"00011011", B"00100010", B"01001000",
 B"00100111", B"11101111", B"11100011", B"00110001", B"00101110",
 B"11011010", B"11101000", B"00111110", B"11011011", B"11101011",
 B"11111010", B"11000110", B"01000011", B"11101100", B"00111010",
 B"00011011", B"11101011", B"00010010", B"00001000", B"11011101",
 B"00100100", B"00010101", B"11001000", B"00010000", B"00011101",
 B"11010000", B"00011010", B"00001011", B"11010111", B"11100101",
 B"00100101", B"11100010", B"00011011", B"00000101", B"11100100",
 B"11110000", B"00011001", B"00011001", B"11100111", B"11010110",
 B"00010010", B"00111001", B"11111001", B"11010101", B"11001100",
 B"11101001", B"11111001", B"00101000", B"11011010", B"11000001",
 B"11011001", B"11101100", B"01000100", B"11010010", B"00001111",
 B"11010010", B"11100000", B"11011110", B"00100101", B"00100100",
 B"11101011", B"00101100", B"11010011", B"00111100", B"00111011",
 B"00110001", B"11101101", B"00100100", B"11100001", B"00010100",
 B"11010000", B"11101100", B"00001100", B"00011000", B"11010100",
 B"11011010", B"11100010", B"11111110", B"11000111", B"00010110",
 B"11101011", B"11100110", B"00011000", B"11101001", B"11110011",
 B"11110001", B"11101011", B"00000010", B"00110001", B"00101000",
 B"11111100", B"11110110", B"11110011", B"11100100", B"10111100",
 B"11110111", B"11001100", B"11010011", B"11010111", B"11111010",
 B"00011000", B"11110100", B"00100110", B"11001111", B"11110010",
 B"11011101", B"11010001", B"00100101", B"00101010", B"00011111",
 B"00101110", B"00001001", B"00011010", B"11110110", B"00110110",
 B"00001001", B"11011111", B"11010110", B"00011101", B"11011011",
 B"00100110", B"11111010", B"00001111", B"11110101", B"11111111",
 B"00100101", B"00011111", B"00010101", B"00011011", B"11011000",
 B"11101010", B"00001000", B"00101011", B"11100010", B"11101010",
 B"00110100", B"11010111", B"00101001", B"11100000", B"11010011",
 B"11011110", B"00110001", B"00010000", B"11011000", B"00110111",
 B"11011101", B"00101001", B"11101101", B"11110010", B"00110010",
 B"00101111", B"00100110", B"00010100", B"00101111", B"00100000",
 B"00011010", B"11101111", B"11111111", B"00100101", B"00011010",
 B"00010011", B"00111100", B"00000001", B"00100000", B"00101110",
 B"00100100", B"00100011", B"00110001", B"00101101", B"00100101",
 B"11100011", B"00010011", B"11010000", B"11111010", B"11010001",
 B"00111100", B"11011000", B"11101110", B"00011101", B"11100101",
 B"11110111", B"11001100", B"11011111", B"11010111", B"10111100",
 B"11001100", B"11010100", B"00000010", B"00001101", B"00010110",
 B"00100111", B"00010110", B"00110010", B"11100111", B"00011001",
 B"11111111", B"11101010", B"11000000", B"00111001", B"00100000",
 B"11011011", B"00110010", B"00011100", B"11010011", B"00100011",
 B"00011011", B"11011110", B"11010111", B"11100111", B"00101110",
 B"00101001", B"00010111", B"00101001", B"11010010", B"00001011",
 B"00010110", B"11010010", B"00101010", B"00101010", B"11011001",
 B"00011001", B"00100000", B"11010100", B"00010101", B"00011110",
 B"00110111", B"00000100", B"00100001", B"11100001", B"00010100",
 B"11101000", B"00101011", B"00100100", B"00101001", B"00010111",
 B"00011110", B"00110001", B"00111100", B"00011111", B"11010110",
 B"00001100", B"11101011", B"00010000", B"11100011", B"11011011",
 B"00010110", B"00010111", B"11101001", B"00100101", B"00100010",
 B"11001100", B"11011101", B"11111000", B"11010011", B"11011000",
 B"11100001", B"00011001", B"11011110", B"11010110", B"11010111",
 B"00111101", B"00010100", B"11100000", B"00001101", B"11011111",
 B"00010110", B"11101011", B"11011100", B"10111100", B"00001011",
 B"00100100", B"11110011", B"11101101", B"00011001", B"11110010",
 B"00100011", B"11101101", B"11011110", B"00100010", B"11011000",
 B"11000111", B"00011001", B"00100010", B"00100001", B"00100000",
 B"11011000", B"11010000", B"00000110", B"00010001", B"11101101",
 B"00101101", B"11101111", B"11101001", B"00010001", B"00011101",
 B"00100011", B"00101011", B"11010000", B"00011010", B"11111101",
 B"11100110", B"11010011", B"00100000", B"11101100", B"11101110",
 B"00011001", B"11011100", B"00101010", B"11100101", B"11010110",
 B"00011001", B"11110111", B"11001110", B"11010101", B"11100111",
 B"00100011", B"00000000", B"00101110", B"00010011", B"11100011",
 B"00011111", B"00011001", B"00010110", B"11101000", B"00001011",
 B"11110010", B"00010110", B"00010011", B"11011111", B"00001011",
 B"11100011", B"11010111", B"01001010", B"11010000", B"00010010",
 B"00011111", B"11100111", B"00110111", B"11111001", B"11100101",
 B"11000100", B"00101100", B"00101100", B"00100000", B"00010111",
 B"11101100", B"00000011", B"00000111", B"11100110", B"11101011",
 B"00110100", B"11011011", B"11011100", B"00001100", B"11010100",
 B"00111010", B"11100001", B"11011011", B"00010100", B"00000111",
 B"11011000", B"11110011", B"11101001", B"11101100", B"00001000",
 B"11110101", B"00100110", B"11101100", B"11011000", B"11010011",
 B"00001000", B"00101000", B"11110001", B"00100110", B"11101100",
 B"11100011", B"00101001", B"11101010", B"11100011", B"11100101",
 B"00100010", B"01001010", B"11001100", B"00101000", B"11100111",
 B"10111110", B"00001111", B"00000001", B"11100100", B"11111010",
 B"11001010", B"00000100", B"11101000", B"00010101", B"11011010",
 B"11100101", B"11010010", B"00100111", B"00101001", B"11011010",
 B"00100000", B"11111001", B"00000111", B"11100001", B"11010100",
 B"00011110", B"00011011", B"11010011", B"00010001", B"00100110",
 B"11100100", B"11011100", B"11100100", B"11101111", B"11011010",
 B"00101110", B"00111101", B"00011000", B"11101110", B"00100101",
 B"11010101", B"00011110", B"11100000", B"00011111", B"00010100",
 B"00011111", B"11001100", B"00100011", B"11011101", B"00010101",
 B"11100100", B"11100101", B"00010101", B"00010001", B"00001101",
 B"11011100", B"00011111", B"11001010", B"00011111", B"00011101",
 B"11001111", B"00111100", B"00010111", B"11100010", B"00010111",
 B"00111011", B"11100101", B"11010110", B"00011010", B"11001111",
 B"00110111", B"11100001", B"11101101", B"00010110", B"01000000",
 B"11011110", B"11100010", B"11100010", B"11011011", B"00001010",
 B"00001101", B"00110011", B"00110010", B"11100000", B"11101000",
 B"01000110", B"00100010", B"00101011", B"00010110", B"11001000",
 B"11011100", B"11100011", B"00101111", B"00101010", B"00011110",
 B"11100011", B"00100111", B"11011111", B"00010000", B"00110011",
 B"11100100", B"00010111", B"11010111", B"11011010", B"11110011",
 B"00101000", B"00011100", B"11011101", B"00001010", B"11100101",
 B"00100000", B"11110110", B"11110100", B"00101011", B"00010111",
 B"00100000", B"00101111", B"11000110", B"11100010", B"00010111",
 B"00011011", B"11100001", B"11101101", B"00101110", B"00010111",
 B"11011000", B"00010111", B"00100101", B"11100001", B"11101010",
 B"00100111", B"11110110", B"00101011", B"11101100", B"00100000",
 B"11111101", B"11010001", B"00110010", B"00010101", B"11001000",
 B"00100000", B"11100001", B"00100111", B"11101010", B"11100100",
 B"00110100", B"00100010", B"00011101", B"11100011", B"11101000",
 B"00101101", B"11100011", B"11011010", B"11010000", B"11100011",
 B"00001110", B"11110011", B"00101000", B"11100111", B"11011001",
 B"11101111", B"00011110", B"00101011", B"00011111", B"00010001",
 B"00011010", B"00011111", B"00011011", B"01000001", B"00011111",
 B"00011011", B"00001100", B"00010101", B"11000010", B"11100011",
 B"00010111", B"00100101", B"11110111", B"11100000", B"00001100",
 B"00010011", B"11111001", B"11100101", B"00011100", B"00010100",
 B"11101010", B"10111100", B"00100010", B"11000011", B"11101010",
 B"00011011", B"11011010", B"11100000", B"11011000", B"11100111",
 B"00000001", B"00101001", B"11101011", B"11011000", B"00010010",
 B"00111001", B"11010000", B"10111111", B"11001101", B"11101011",
 B"00100101", B"00011000", B"00011010", B"00100001", B"11001100",
 B"11010001", B"11110010", B"11010111", B"11110000", B"11101101",
 B"11111001", B"00100110", B"00011110", B"00110000", B"01000011",
 B"00110101", B"00011011", B"11100000", B"01010010", B"11010101",
 B"00101010", B"10111011", B"11101011", B"11110000", B"00010001",
 B"11010110", B"00011111", B"11001100", B"11010010", B"00010000",
 B"11011010", B"00010010", B"11010011", B"11100110", B"11010111",
 B"00101001", B"00010111", B"11010110", B"11100000", B"11101100",
 B"11001011", B"11100100", B"00010011", B"00001001", B"00000101",
 B"00000111", B"11001101", B"11001001", B"00011101", B"00001010",
 B"00011011", B"00101101", B"11011111", B"11101111", B"00000011",
 B"00011101", B"00010000", B"00101000", B"11011100", B"00100111",
 B"11001111", B"00011110", B"11110101", B"00110011", B"11011100",
 B"00000100", B"00011011", B"11011011", B"11101011", B"00011101",
 B"11001110", B"11001000", B"00001110", B"00011110", B"00011111",
 B"00001011", B"11100110", B"00000011", B"00011100", B"00011100",
 B"11010101", B"00100010", B"00011111", B"11100000", B"11110000",
 B"00100000", B"11101001", B"11100011", B"00100010", B"00010000",
 B"00100100", B"00010111", B"11100001", B"11111010", B"00101001",
 B"00011100", B"00100001", B"11011111", B"00100111", B"11010000",
 B"00110000", B"11110111", B"11100011", B"11001100", B"00001000",
 B"11101000", B"00100101", B"11010000", B"00000111", B"00001001",
 B"00100101", B"11101111", B"11101010", B"11101011", B"11100010",
 B"00010110", B"11010010", B"00100001", B"00011010", B"00100110",
 B"00011011", B"11010010", B"00001010", B"11010000", B"00010000",
 B"11011000", B"11100101", B"11011100", B"11101110", B"00101101",
 B"00110010", B"11111101", B"00100011", B"11101001", B"11101011",
 B"00100111", B"11101010", B"00001110", B"11011100", B"11100000",
 B"00110011", B"00101111", B"00001011", B"00011000", B"11001111",
 B"00011001", B"00100101", B"11001111", B"11101001", B"00100110",
 B"11110101", B"11011101", B"11101110", B"11000111", B"00000010",
 B"00101100", B"00100101", B"00100111", B"00111111", B"11010111",
 B"00011001", B"11011110", B"11100000", B"11010111", B"00101100",
 B"00100111", B"11110111", B"00011110", B"11111010", B"11101111",
 B"11110001", B"00100000", B"00011101", B"11011010", B"11111001",
 B"11100110", B"11010101", B"00011100", B"00100001", B"11101010",
 B"00011011", B"11011111", B"00100110", B"00010110", B"00101001",
 B"11110100", B"01000010", B"11101000", B"00101000", B"11111110",
 B"00010111", B"00011001", B"00001011", B"11101100", B"00011100",
 B"11111000", B"00010000", B"11010110", B"11100011", B"00010011",
 B"00110111", B"00011100", B"11111101", B"00110100", B"11011111",
 B"00111111", B"11101001", B"00100001", B"00010000", B"00100001",
 B"11100110", B"00100110", B"00001011", B"00011001", B"11010010",
 B"00011101", B"00110001", B"00010100", B"11111010", B"00110001",
 B"11110111", B"00111010", B"11101000", B"00010001", B"11100101",
 B"11100110", B"11011111", B"00100011", B"00000001", B"11000101",
 B"00011011", B"11101000", B"01000000", B"11101111", B"11100100",
 B"11010000", B"00000110", B"00100110", B"11010100", B"00101011",
 B"00011000", B"00011101", B"11011111", B"00001100", B"11001011",
 B"00001011", B"11110010", B"00110010", B"11010010", B"11100110",
 B"11011100", B"00010110", B"00101010", B"11011110", B"00110001",
 B"00011110", B"11110100", B"11011010", B"00011100", B"00100001",
 B"11001001", B"11110010", B"00000111", B"00101010", B"00111000",
 B"11110000", B"00101010", B"11000101", B"00101001", B"11110101",
 B"11011100", B"11011010", B"11000010", B"00100100", B"00111100",
 B"11010110", B"00111111", B"11010101", B"11100111", B"11111000",
 B"11110000", B"11100011", B"11111001", B"00110011", B"00010110",
 B"00101001", B"00001001", B"11001010", B"11100111", B"11010111",
 B"11110010", B"00101110", B"11010011", B"00001011", B"00010000",
 B"00100000", B"11010000", B"00001101", B"00001001", B"11100110",
 B"11010000", B"00100100", B"00001110", B"11100101", B"00110101",
 B"11001011", B"11010110", B"11101101", B"00000100", B"00100011",
 B"00111001", B"11010101", B"10111001", B"00010010", B"11011010",
 B"11101001", B"11011111", B"11101111", B"00110100", B"00011000",
 B"00011011", B"00110100", B"00101001", B"00010001", B"00011011",
 B"00000111", B"11100011", B"11110000", B"11110011", B"00011101",
 B"00011011", B"11100111", B"00011101", B"11100011", B"00101111",
 B"00011100", B"00100110", B"00111100", B"00101010", B"00010000",
 B"00100111", B"00100011", B"00010101", B"11100010", B"11100111",
 B"11101011", B"11010111", B"11100111", B"11011000", B"11100000",
 B"11011000", B"00011110", B"11100011", B"11101010", B"11111101",
 B"00101011", B"00101011", B"11110000", B"00001100", B"11011110",
 B"00001100", B"11110110", B"11011001", B"11010110", B"00000100",
 B"00010100", B"00011010", B"00011111", B"00110111", B"11010110",
 B"00100010", B"11111010", B"01000110", B"11111100", B"00101010",
 B"00011001", B"00100100", B"11001111", B"11111001", B"11001001",
 B"01000011", B"11100001", B"11100100", B"11011111", B"11101101",
 B"11001000", B"00010010", B"00101010", B"00010001", B"00111010",
 B"11011010", B"11110010", B"00010101", B"00011001", B"11110100",
 B"00110111", B"11101111", B"11101011", B"11010011", B"11011111",
 B"11110111", B"00010100", B"00101011", B"11110001", B"00100011",
 B"11011011", B"00010100", B"00101011", B"00100011", B"00110010",
 B"00111101", B"00101110", B"01000011", B"00001111", B"00101110",
 B"11011011", B"00101001", B"11000101", B"11110101", B"11001101",
 B"00100111", B"00011001", B"11010000", B"00100111", B"11010010",
 B"11011011", B"11010101", B"00111011", B"00101001", B"11100100",
 B"11111110", B"00100010", B"11101100", B"11101001", B"11110111",
 B"00001110", B"01001001", B"11110100", B"00000010", B"00110100",
 B"00100000", B"00010110", B"00010101", B"00101101", B"00100001",
 B"00100101", B"00101111", B"11101110", B"11001111", B"00010101",
 B"11100101", B"11011111", B"11110101", B"11100001", B"00010001",
 B"11011011", B"11011111", B"11001101", B"11010111", B"01001110",
 B"11100110", B"00101110", B"00011001", B"11100110", B"11110001",
 B"11011101", B"11000110", B"00010111", B"11010110", B"00010111",
 B"11100101", B"10110001", B"11100101", B"00011010", B"00100010",
 B"11000000", B"00011100", B"11101011", B"00100011", B"00101001",
 B"11110110", B"11101011", B"00011101", B"00010001", B"11101000",
 B"11100100", B"00000111", B"11110101", B"00010101", B"00100110",
 B"01000000", B"00011001", B"00010110", B"00010111", B"11001001",
 B"00000100", B"00011000", B"00100101", B"00111001", B"00000000",
 B"11001110", B"11010111", B"00011110", B"11011100", B"11001100",
 B"00110011", B"11110011", B"11100110", B"11100000", B"11010101",
 B"00100100", B"00011100", B"00011010", B"00101111", B"00010100",
 B"00001111", B"00100111", B"00011000", B"11011011", B"00011010",
 B"00011000", B"00101010", B"10110010", B"00100110", B"11011011",
 B"00111011", B"00100000", B"00010010", B"11100100", B"00100111",
 B"00110111", B"11101100", B"11010101", B"00100101", B"00011010",
 B"11101011", B"00100111", B"00010000", B"11011010", B"00110010",
 B"00001111", B"11101110", B"11010101", B"11101001", B"00011000",
 B"11110010", B"00101011", B"11011101", B"11010011", B"11111101",
 B"00001011", B"00010101", B"00000100", B"00111001", B"00101100",
 B"00001111", B"00110010", B"00101110", B"00101100", B"00010110",
 B"00101100", B"00011110", B"00011110", B"00011001", B"00011100",
 B"00101101", B"00011101", B"00001111", B"00000011", B"11010111",
 B"00000100", B"11001100", B"00010011", B"11101110", B"00100111",
 B"11010110", B"00100101", B"00000101", B"11100010", B"00101000",
 B"00011110", B"11101101", B"11100111", B"11101100", B"00010111",
 B"11011110", B"00110011", B"11011000", B"00000110", B"00110100",
 B"00011111", B"00100011", B"11111100", B"11010000", B"00011001",
 B"00100101", B"11101001", B"11010110", B"11001111", B"00110010",
 B"00100001", B"11011000", B"11101001", B"11101010", B"11011111",
 B"11000110", B"00011111", B"11100000", B"11100100", B"00001010",
 B"11100101", B"11100111", B"11110011", B"11010001", B"11011101",
 B"00110101", B"00100111", B"11111011", B"11000101", B"11011101",
 B"11100011", B"11101010", B"01000010", B"00101010", B"11110000",
 B"00001101", B"00010111", B"00100110", B"00101100", B"00101010",
 B"00100101", B"00100100", B"00010111", B"00011101", B"00101100",
 B"00110001", B"00011001", B"00110010", B"00011001", B"00100110",
 B"00010111", B"11101111", B"00101010", B"11110110", B"00110111",
 B"11100000", B"11011111", B"00000011", B"11100110", B"11011000",
 B"11110000", B"00110110", B"00011110", B"11100100", B"11011111",
 B"00011010", B"00001110", B"00010011", B"10111110", B"00010010",
 B"11010110", B"00010111", B"11010011", B"00010100", B"00010000",
 B"11110011", B"11011011", B"11011101", B"11010000", B"11101101",
 B"00011000", B"11111000", B"00010011", B"00010100", B"00100100",
 B"00011010", B"00010110", B"00100101", B"11100000", B"00100000",
 B"00010000", B"00101101", B"11111011", B"00100100", B"11000010",
 B"00101111", B"11101100", B"11101110", B"00011100", B"11101111",
 B"00011011", B"11010111", B"11110010", B"00011111", B"00011010",
 B"11111110", B"11100100", B"11011100", B"11011101", B"00011101",
 B"11011101", B"00010101", B"00100100", B"11101010", B"11110110",
 B"11111100", B"11100001", B"00000100", B"11111010", B"11101011",
 B"00110111", B"11011110", B"00100001", B"00001111", B"11000110",
 B"00100101", B"01001011", B"11111001", B"11101001", B"00011010",
 B"11011110", B"11101111", B"11101010", B"00110011", B"00100011",
 B"11001110", B"00101001", B"00110000", B"11111010", B"00100101",
 B"00011100", B"11110001", B"11101000", B"00011011", B"00100110",
 B"00101011", B"00010011", B"00111001", B"00000011", B"01000010",
 B"00010001", B"00011111", B"01000100", B"11001001", B"00100111",
 B"00101011", B"11010100", B"00010110", B"00001011", B"10111011",
 B"11110111", B"00011000", B"11010100", B"00101010", B"11100100",
 B"11110101", B"00110110", B"00011010", B"11000000", B"11001000",
 B"00010001", B"11100100", B"00001110", B"11001000", B"11100100",
 B"00110010", B"11100010", B"00011000", B"11110110", B"11110100",
 B"11110010", B"00011000", B"00100011", B"11101101", B"11110011",
 B"10111000", B"00011001", B"00010111", B"00011010", B"00100101",
 B"11000100", B"11010110", B"00001111", B"11010100", B"11010101",
 B"11110001", B"11010100", B"00011101", B"11000111", B"00100110",
 B"11011011", B"11001010", B"11110010", B"11011101", B"00101110",
 B"00011110", B"00001111", B"00001101", B"00100011", B"11000100",
 B"11100010", B"00010001", B"11110100", B"11011100", B"11100101",
 B"11011000", B"01000001", B"00010111", B"11010011", B"11001101",
 B"00100000", B"00011110", B"11110011", B"11101000", B"00101010",
 B"00000101", B"00011111", B"11010011", B"00101100", B"11010000",
 B"00001110", B"11011101", B"00010100", B"11010111", B"00010101",
 B"00100011", B"11001111", B"00011101", B"00010101", B"11001101",
 B"00000111", B"00011011", B"00100100", B"11011101", B"00110010",
 B"11110000", B"00011000", B"11001001", B"11100001", B"00100000",
 B"11110100", B"00110010", B"11000001", B"11101111", B"00010010",
 B"00000110", B"11010010", B"00101010", B"11011011", B"11101100",
 B"11011000", B"00110001", B"00100100", B"11100100", B"00011011",
 B"00001001", B"11001011", B"00001001", B"11000111", B"11110111",
 B"11100111", B"11100000", B"11011101", B"11011110", B"11101101",
 B"11000111", B"00101010", B"00000110", B"00101000", B"00101101",
 B"00001001", B"00111010", B"11101001", B"00010101", B"11101010",
 B"11100011", B"00100011", B"00011101", B"11011001", B"11001010",
 B"11010101", B"00110100", B"00100100", B"11100010", B"00101010",
 B"11110011", B"00001111", B"00110011", B"11001111", B"00101100",
 B"00011101", B"11101000", B"11010101", B"00101010", B"11101111",
 B"00010011", B"00101000", B"00101100", B"11100101", B"00101111",
 B"11001000", B"00010000", B"00011101", B"11011010", B"00011001",
 B"00101110", B"11000111", B"00100100", B"00010111", B"11110001",
 B"00011111", B"01000001", B"11011000", B"00110001", B"00110100",
 B"11101010", B"11010111", B"00000011", B"10111100", B"00111111",
 B"11101010", B"00110011", B"11100010", B"11001001", B"00101001",
 B"00110001", B"11001000", B"00100001", B"11110110", B"00010110",
 B"11001111", B"11001100", B"00011011", B"00010000", B"11011010",
 B"00010111", B"11110110", B"00010011", B"11010101", B"11010100",
 B"00110001", B"00011000", B"00011110", B"00010100", B"00100110",
 B"11011110", B"00000011", B"11100101", B"00011000", B"11010111",
 B"00000101", B"00111011", B"11011001", B"00111101", B"11111010",
 B"11100110", B"00111110", B"00101010", B"00110011", B"00101001",
 B"00011011", B"00101000", B"00011001", B"00011100", B"00001111",
 B"00101110", B"11010011", B"00101011", B"11101100", B"00111101",
 B"11111100", B"00001000", B"00101111", B"00001111", B"00010110",
 B"10111100", B"00010010", B"11011110", B"11100001", B"11000011",
 B"00110001", B"00101010", B"11010110", B"01000110", B"11100100",
 B"11010000", B"11010101", B"00100110", B"00001101", B"11011011",
 B"00101101", B"01001100", B"00111011", B"00101000", B"00010000",
 B"00110100", B"00100000", B"00011100", B"00100101", B"11100111",
 B"00101010", B"00100100", B"11010001", B"00001010", B"00110000",
 B"11100111", B"11010011", B"00001101", B"00001101", B"00010000",
 B"11110111", B"00101010", B"11100000", B"00100100", B"11101100",
 B"11100010", B"11011011", B"11101000", B"00101100", B"00101110",
 B"00010110", B"00011111", B"00110011", B"11011111", B"00100000",
 B"00101111", B"11110001", B"00100010", B"00011001", B"11010110",
 B"11110101", B"00011110", B"11110001", B"00011011", B"11100110",
 B"11001001", B"00110001", B"11101110", B"11011101", B"11010100",
 B"10111101", B"11000011", B"00100000", B"00111101", B"00010010",
 B"00101010", B"11011111", B"00010110", B"00010001", B"00101010",
 B"11110010", B"00011000", B"11100100", B"00101011", B"11011000",
 B"11001100", B"11010010", B"00110000", B"00110000", B"11100001",
 B"00110100", B"11100101", B"00011001", B"00001010", B"11000101",
 B"11110110", B"11100011", B"00101110", B"00000111", B"00010000",
 B"11011100", B"10111001", B"11010001", B"00000110", B"00011100",
 B"11011101", B"00110001", B"11011011", B"11000000", B"00110010",
 B"11001110", B"11111101", B"11001000", B"00101000", B"00110010",
 B"11100011", B"00101000", B"00111011", B"00000010", B"00010010",
 B"01000010", B"00010101", B"00011010", B"00010000", B"11010100",
 B"11011011", B"00110100", B"00011110", B"00100110", B"00011000",
 B"11110010", B"11001110", B"00001111", B"00101110", B"11010100",
 B"11001000", B"00110100", B"00010111", B"11011010", B"11011010",
 B"00100000", B"00011001", B"00100111", B"00100100", B"00110001",
 B"00100000", B"00001001", B"00010100", B"11001111", B"00011100",
 B"11111001", B"11011101", B"11010110", B"00100010", B"01000100",
 B"11101101", B"11010100", B"11011101", B"00010111", B"00100111",
 B"00110100", B"00000010", B"11010101", B"11010111", B"00100000",
 B"00010110", B"11011110", B"00101001", B"00101111", B"11011110",
 B"11010110", B"00010111", B"11111100", B"00100000", B"00101111",
 B"00110001", B"11101010", B"00011001", B"11101100", B"00011001",
 B"11010111", B"00011100", B"11011101", B"11100011", B"11011100",
 B"00010011", B"00011110", B"11101011", B"00101010", B"11100111",
 B"11101101", B"00011101", B"11000101", B"11101100", B"11001100",
 B"11001101", B"11000101", B"00011010", B"00011000", B"00101111",
 B"11100111", B"00100011", B"11001000", B"00110101", B"11110100",
 B"11010110", B"11000001", B"11100011", B"00101011", B"00010100",
 B"00010110", B"00100101", B"11100111", B"00001010", B"11111011",
 B"00110001", B"11010010", B"00100100", B"11110011", B"00100010",
 B"00100101", B"11100011", B"11100000", B"00011101", B"11011100",
 B"11100101", B"11110010", B"11100000", B"11100100", B"11011000",
 B"00011000", B"00010101", B"01000011", B"00100001", B"11011101",
 B"11110110", B"11101110", B"00010100", B"00001010", B"11001110",
 B"11100100", B"11011000", B"11111010", B"11010110", B"11011100",
 B"10111011", B"00111011", B"11010100", B"00110010", B"11001100",
 B"11011100", B"00111000", B"11011110", B"00011101", B"00100011",
 B"11011111", B"11100010", B"11101000", B"11010111", B"11011101",
 B"00001110", B"00100100", B"11011111", B"00110000", B"00011111",
 B"11011000", B"11001010", B"00111010", B"00011111", B"11101000",
 B"00011111", B"11111111", B"11011010", B"00110011", B"01000100",
 B"11100111", B"00001001", B"11101100", B"00011000", B"11011001",
 B"11011111", B"11100111", B"00010011", B"00101001", B"01000100",
 B"11101001", B"00100110", B"11010001", B"11011101", B"11110000",
 B"00010110", B"00010111", B"11010100", B"00110101", B"11101101",
 B"00001101", B"11101000", B"11100101", B"00111001", B"00000110",
 B"00100010", B"00010110", B"00101101", B"00110001", B"00010010",
 B"00010110", B"00000101", B"00100000", B"11101111", B"00001000",
 B"00111001", B"00010101", B"00001100", B"00010011", B"11111000",
 B"00011111", B"11110000", B"00010011", B"11111000", B"00110000",
 B"11101011", B"11101000", B"11111101", B"00100011", B"11101101",
 B"11100011", B"00010110", B"00110111", B"00101011", B"00001101",
 B"11010101", B"11100110", B"00110001", B"11101000", B"11110011",
 B"00101011", B"11101101", B"11100010", B"11011101", B"11011111",
 B"00101000", B"11101110", B"11010101", B"00101101", B"11101111",
 B"11110000", B"11010000", B"11010111", B"11010101", B"11101101",
 B"00011010", B"00011011", B"00011001", B"00011101", B"11011111",
 B"11001011", B"00100111", B"00111100", B"11100001", B"11011000",
 B"11111100", B"00110011", B"11010110", B"11100000", B"00101011",
 B"00001000", B"11010011", B"00001010", B"00011000", B"11101000",
 B"11000010", B"00100001", B"00011001", B"00101011", B"00100001",
 B"11111110", B"00100110", B"00010100", B"00111000", B"00011110",
 B"00011010", B"11001010", B"01010011", B"00101001", B"11011010",
 B"00100001", B"00011010", B"11101010", B"00001110", B"00010101",
 B"11001111", B"00000000", B"00110001", B"11101011", B"11110100",
 B"00110111", B"11100100", B"00001011", B"11100110", B"00100100",
 B"11011011", B"11001100", B"00101010", B"00101100", B"11110101",
 B"00100010", B"11100001", B"00110010", B"11101100", B"10111111",
 B"00001100", B"00101001", B"00001011", B"11010111", B"00111010",
 B"11010110", B"11100101", B"11101001", B"00011000", B"00101100",
 B"00100111", B"11010111", B"11100100", B"00101101", B"11100010",
 B"11101101", B"11101011", B"11010111", B"11101101", B"00001100",
 B"00100010", B"00110100", B"11100100", B"00101000", B"11101111",
 B"00010000", B"00111101", B"00011000", B"00100101", B"11100110",
 B"00100011", B"11011010", B"00010100", B"00000000", B"00100101",
 B"11000101", B"00010011", B"00010111", B"11110001", B"01000010",
 B"11110110", B"11011101", B"11010110", B"11010000", B"11101010",
 B"11011011", B"00011101", B"00011011", B"00100000", B"00010100",
 B"00101010", B"00011011", B"10111100", B"11001011", B"00011001",
 B"00110100", B"11110111", B"11110000", B"00001001", B"11101100",
 B"11101110", B"11011111", B"11100110", B"00011010", B"11011011",
 B"00010000", B"11011011", B"00100100", B"00100010", B"11101010",
 B"11010110", B"11000011", B"11110001", B"11110010", B"00100100",
 B"11110001", B"11001100", B"11011101", B"11010011", B"00111110",
 B"11101011", B"00001101", B"00010011", B"11001101", B"11101000",
 B"00100000", B"10110101", B"11011110", B"11001101", B"11010000",
 B"11100000", B"11011111", B"00100000", B"00011110", B"00101011",
 B"00010101", B"11011011", B"11100110", B"11101001", B"00010011",
 B"11011010", B"00100001", B"11110111", B"11111111", B"00101001",
 B"00011001", B"11100101", B"00001111", B"00011000", B"11010010",
 B"11010110", B"11110011", B"11100110", B"10111000", B"00010110",
 B"00110000", B"11100011", B"11100000", B"00100001", B"00010011",
 B"11010111", B"11001110", B"00001111", B"00011000", B"00001111",
 B"00100100", B"00100101", B"00111010", B"00110011", B"00001010",
 B"00011011", B"00110111", B"11100101", B"00011001", B"00001110",
 B"11101001", B"11101011", B"00111101", B"00011000", B"11101101",
 B"11011110", B"00011101", B"11011101", B"11100111", B"11101011",
 B"11110011", B"00001000", B"00001100", B"00100101", B"00110001",
 B"00101001", B"00100010", B"00001000", B"00010100", B"11010101",
 B"11100111", B"00000111", B"00101101", B"00100001", B"00010111",
 B"11100111", B"11010111", B"11011011", B"11101001", B"00101111",
 B"11001110", B"00100101", B"11011001", B"11011000", B"00100011",
 B"00101100", B"10111111", B"00101010", B"00110011", B"11100000",
 B"00101110", B"00011110", B"11100011", B"00101100", B"00010100",
 B"11100010", B"11111101", B"00101011", B"11011001", B"11100000",
 B"00101101", B"11011101", B"11110000", B"11001101", B"00100000",
 B"00100101", B"11100010", B"00101010", B"11000000", B"00001010",
 B"00110001", B"11100111", B"11100000", B"00001001", B"00100000",
 B"11110000", B"11111011", B"00100100", B"00110011", B"00100010",
 B"11110111", B"00101101", B"11111100", B"00110000", B"11110101",
 B"10111101", B"00010100", B"11011011", B"11100100", B"11011000",
 B"00100110", B"00110111", B"11100011", B"00101111", B"00110101",
 B"00110000", B"00010000", B"00000011", B"00011011", B"00100010",
 B"00000101", B"11010110", B"00010001", B"11110100", B"00101111",
 B"11111010", B"11110001", B"00011111", B"00110011", B"00100001",
 B"00011001", B"11011100", B"11100010", B"00010011", B"00010111",
 B"11101001", B"11011101", B"00100001", B"00110101", B"11111011",
 B"11001100", B"00010100", B"00010010", B"00000010", B"11001000",
 B"00101110", B"11101110", B"11001110", B"11100000", B"11111000",
 B"00011100", B"11011010", B"00110111", B"00101101", B"11011101",
 B"00110101", B"00100001", B"11010010", B"00110110", B"00101011",
 B"11110000", B"00101111", B"00001111", B"00001101", B"11010111",
 B"00100011", B"11111010", B"00001110", B"11100001", B"11010000",
 B"11100111", B"00010100", B"00010110", B"00011110", B"00100001",
 B"11011101", B"11010111", B"11010110", B"00101011", B"00011111",
 B"00001101", B"11000110", B"00000000", B"11001100", B"00011000",
 B"11101110", B"11011100", B"00001100", B"11100100", B"11111100",
 B"11011001", B"11001101", B"00110110", B"00011001", B"11100010",
 B"00010001", B"00100011", B"11100100", B"00100001", B"00011001",
 B"11011011", B"11111000", B"11101111", B"00111111", B"11100111",
 B"00110001", B"11100101", B"11110001", B"00100010", B"00000111",
 B"00010110", B"11100101", B"00100010", B"00011111", B"11011000",
 B"11100001", B"00101011", B"11101111", B"00001111", B"11100110",
 B"11100010", B"11100011", B"00101010", B"00010111", B"11001110",
 B"11101011", B"00001101", B"11110111", B"00010010", B"11001010",
 B"11100111", B"00010110", B"11111100", B"11101000", B"00010111",
 B"11011111", B"11010101", B"10111100", B"00001010", B"00101110",
 B"11101101", B"00010111", B"00101100", B"11011101", B"11001111",
 B"00100101", B"00010010", B"00000010", B"11100011", B"11011101",
 B"00000001", B"00011100", B"00011000", B"11101110", B"00100000",
 B"11100100", B"00101100", B"11110011", B"00110110", B"00011000",
 B"00100110", B"11101001", B"00110111", B"11010011", B"00001001",
 B"00101111", B"00111110", B"11011001", B"00110011", B"00000011",
 B"11110111", B"11100100", B"00100110", B"11100010", B"00011111",
 B"11100000", B"00001001", B"11100101", B"11101011", B"00110111",
 B"00110010", B"00101110", B"00110001", B"11001100", B"00100110",
 B"00100111", B"11100011", B"11011111", B"00001111", B"00010011",
 B"11110010", B"11101101", B"00110111", B"11110101", B"11100000",
 B"11010000", B"11110110", B"11101011", B"11011011", B"00001010",
 B"00111010", B"00011011", B"00110011", B"11101101", B"11100100",
 B"11011000", B"11100111", B"11100000", B"00101010", B"00001110",
 B"11001101", B"00100100", B"11011111", B"00010011", B"00100010",
 B"11001011", B"00011010", B"00011100", B"11000101", B"11100110",
 B"00101000", B"00011001", B"11001011", B"11011011", B"00011110",
 B"11101011", B"11110010", B"11010010", B"11101011", B"00010000",
 B"00100011", B"00011100", B"11001000", B"00001010", B"11100101",
 B"01000000", B"11010110", B"00000010", B"11010110", B"11101111",
 B"11010100", B"11100000", B"00101011", B"11101100", B"00100110",
 B"11001100", B"11001011", B"00000111", B"11101011", B"00100111",
 B"11101110", B"11100000", B"00010100", B"11010110", B"11110000",
 B"00100001", B"11010001", B"00111111", B"11101110", B"11101000",
 B"00001010", B"11100101", B"11001110", B"11010101", B"11100111",
 B"00100011", B"00101100", B"00100000", B"00001011", B"00101110",
 B"00011111", B"11110110", B"00011011", B"00010001", B"11100001",
 B"11011010", B"00010111", B"00011111", B"00010000", B"00011111",
 B"11011011", B"00001100", B"11101100", B"00100111", B"11000011",
 B"00100010", B"00110100", B"11101010", B"11001110", B"00001011",
 B"00110011", B"11110000", B"11000010", B"00110101", B"11010100",
 B"11010010", B"00100100", B"11011000", B"11001001", B"11100101",
 B"11111000", B"00011101", B"11111001", B"00010100", B"00101101",
 B"11011101", B"00110011", B"00011111", B"11011110", B"00010010",
 B"11011010", B"00010011", B"11001110", B"11011011", B"11000111",
 B"00010001", B"00011001", B"10111110", B"00101100", B"00010110",
 B"11101101", B"11111100", B"11001110", B"11100000", B"11101101",
 B"00001011", B"00100000", B"11100011", B"11100011", B"00101110",
 B"00011000", B"11010100", B"11101010", B"00011011", B"00110100",
 B"00101100", B"00100010", B"11111111", B"00010000", B"00011010",
 B"11111001", B"00001111", B"11101011", B"01000101", B"11101001",
 B"11100000", B"11100011", B"00100001", B"00100000", B"11010001",
 B"11100010", B"11010011", B"11100100", B"00101000", B"00101111",
 B"00011101", B"00011101", B"00011001", B"00100011", B"11000111",
 B"00101110", B"00001110", B"11101111", B"11100001", B"01000011",
 B"11100100", B"11100001", B"11011110", B"00010000", B"00001010",
 B"11010111", B"00010100", B"11101000", B"11100011", B"00111001",
 B"11011101", B"00101001", B"11100100", B"11100101", B"00101110",
 B"00100000", B"11100011", B"11010011", B"11100000", B"11101101",
 B"00001111", B"00101011", B"00101000", B"00110011", B"00001100",
 B"00001111", B"11101111", B"11010000", B"00011101", B"00010001",
 B"11010010", B"11100101", B"11101110", B"11010101", B"00100110",
 B"11100010", B"00111010", B"11011011", B"11100110", B"00011000",
 B"00000001", B"00110110", B"11111001", B"11011100", B"00001100",
 B"00101100", B"11000000", B"10110111", B"00011001", B"00001101",
 B"00101111", B"00100010", B"00100111", B"00011001", B"00010110",
 B"00110011", B"00100010", B"11110000", B"00100010", B"11111101",
 B"11010111", B"11000001", B"00100000", B"00010100", B"00011101",
 B"00100010", B"11110111", B"11100011", B"00100100", B"00011100",
 B"11010001", B"11100001", B"00010111", B"11110011", B"00101110",
 B"00101000", B"11010100", B"00011000", B"00100000", B"11100111",
 B"00011000", B"11100111", B"00011001", B"11001111", B"11100101",
 B"00000101", B"00110111", B"00100010", B"00000101", B"11011111",
 B"11111010", B"11001101", B"11111110", B"00011111", B"11100011",
 B"00011100", B"11000011", B"11100001", B"00111110", B"00100000",
 B"00001110", B"11111000", B"11110001", B"11000110", B"00101010",
 B"00001000", B"00101001", B"11101010", B"00001000", B"00000101",
 B"00011001", B"00100010", B"00011001", B"00001010", B"11101100",
 B"00100001", B"00111001", B"11011010", B"11010111", B"00011101",
 B"11101100", B"11010001", B"00110000", B"11101101", B"00101111",
 B"11001010", B"11000011", B"00011011", B"00010100", B"00011000",
 B"11101001", B"00010100", B"00000100", B"11010100", B"11010000",
 B"00011110", B"11100011", B"11000111", B"00011001", B"00101001",
 B"00101000", B"00011001", B"11101000", B"11110111", B"11010110",
 B"11010011", B"11100101", B"00101101", B"00010001", B"11011001",
 B"00001010", B"11100011", B"11010100", B"11101101", B"11110001",
 B"00010111", B"00111110", B"11011110", B"00011110", B"11111010",
 B"00110110", B"00101110", B"11100001", B"11100001", B"00010010",
 B"00011010", B"11101010", B"11011011", B"00100010", B"11001011",
 B"00110010", B"11011101", B"11010111", B"11001011", B"00101110",
 B"00001111", B"11100110", B"00100001", B"00000110", B"11011100",
 B"11100111", B"11011010", B"11001111", B"11010000", B"00011101",
 B"11100010", B"11100001", B"11101001", B"11011110", B"00011010",
 B"11111100", B"00110101", B"00110111", B"00001110", B"00000101",
 B"11110010", B"00111000", B"11101001", B"00110011", B"11011100",
 B"00101001", B"00101110", B"11100000", B"11101011", B"00010110",
 B"00001101", B"11100011", B"11010010", B"11010000", B"00001011",
 B"00010111", B"00010001", B"11011010", B"00100101", B"11100000",
 B"11111111", B"11111100", B"00011100", B"11011111", B"00011011",
 B"00001001", B"11100000", B"11101101", B"00011101", B"00101100",
 B"00111011", B"00011001", B"11001100", B"00010110", B"11011010",
 B"00001101", B"11101111", B"11011111", B"00001110", B"00011000",
 B"00110000", B"11111000", B"00100010", B"11101110", B"11110101",
 B"11100010", B"00101011", B"11001011", B"00011101", B"11100000",
 B"11100010", B"00100101", B"00100101", B"00100011", B"11011011",
 B"11100111", B"00010101", B"11001100", B"11000010", B"11100010",
 B"11101110", B"00011000", B"11100100", B"00100110", B"11111100",
 B"11100101", B"11111010", B"00101110", B"00010001", B"00101101",
 B"00011011", B"11011000", B"00001011", B"00011111", B"11111100",
 B"11011010", B"00101110", B"00101100", B"11010101", B"00010110",
 B"11101110", B"11011110", B"11111001", B"00100011", B"00100100",
 B"00110101", B"00101011", B"11010110", B"00100111", B"00101101",
 B"11010010", B"11001110", B"00101101", B"11101100", B"00110011",
 B"11010101", B"10110001", B"11011101", B"00010100", B"01000011",
 B"11101001", B"11111111", B"11010101", B"11011100", B"11101010",
 B"00100000", B"00000001", B"00010110", B"00110100", B"11011000",
 B"11011111", B"11100000", B"00011100", B"00001110", B"11001000",
 B"00100000", B"11111110", B"00011100", B"11011110", B"00100110",
 B"00001111", B"11110001", B"00010010", B"00011110", B"11101101",
 B"00011000", B"11100011", B"11100011", B"00100010", B"11001100",
 B"11100101", B"11100111", B"11010011", B"11101001", B"00001001",
 B"00010111", B"11001000", B"11011011", B"11001000", B"11010011",
 B"11010101", B"00101101", B"11110100", B"11001110", B"00100111",
 B"11111011", B"11001111", B"11100010", B"11101001", B"00111101",
 B"11111000", B"11100110", B"00000010", B"11011011", B"00110011",
 B"11010010", B"00001011", B"00101100", B"11011100", B"11110011",
 B"11010101", B"11011011", B"00100111", B"11100100", B"00101000",
 B"11010010", B"00011101", B"00101111", B"00100010", B"11001111",
 B"00010010", B"11001111", B"01000111", B"00100011", B"00100000",
 B"00001101", B"11010101", B"00010111", B"11100100", B"00000111",
 B"11011000", B"00000111", B"11010100", B"11101110", B"11100100",
 B"11100110", B"00101100", B"11010000", B"00100100", B"11101000",
 B"11101001", B"00110001", B"11011010", B"00110010", B"11101001",
 B"11010110", B"00100100", B"11111000", B"11001010", B"11101000",
 B"00011000", B"11110101", B"11011111", B"00111110", B"11011011",
 B"11110111", B"00100011", B"11100111", B"11111001", B"11001100",
 B"00011000", B"00101001", B"11110000", B"11010101", B"11100010",
 B"11011010", B"11100011", B"00100101", B"00101100", B"00001000",
 B"00101111", B"00000011", B"00011011", B"11001000", B"00011100",
 B"00010100", B"11101110", B"11111100", B"00101010", B"00010010",
 B"11100010", B"00101011", B"00000110", B"11110111", B"00101100",
 B"00101010", B"00011101", B"11100001", B"11010001", B"00000111",
 B"00010110", B"00100110", B"11101001", B"00000110", B"11010101",
 B"00100111", B"11101001", B"11011111", B"11110011", B"10111010",
 B"00010000", B"11100011", B"00011000", B"00011001", B"00100111",
 B"00000100", B"00010110", B"00100011", B"00011110", B"00010110",
 B"01001101", B"11011110", B"00100110", B"11100001", B"11100110",
 B"11101011", B"00100111", B"00101011", B"11111110", B"00100011",
 B"00101010", B"00101100", B"11100001", B"00100010", B"11010111",
 B"00101110", B"11010101", B"00000011", B"00100001", B"00000010",
 B"00101101", B"00011000", B"11100110", B"11100000", B"00010101",
 B"00101110", B"00101000", B"00011110", B"00011101", B"00001011",
 B"00100011", B"00111111", B"00001011", B"11011101", B"00101000",
 B"11011001", B"11011001", B"11010110", B"00100110", B"00011000",
 B"11001110", B"00010110", B"00010110", B"00011111", B"01000000",
 B"00110001", B"00101011", B"00000101", B"00011010", B"00010110",
 B"11110110", B"00011110", B"11101111", B"11100010", B"11110000",
 B"00101001", B"00100111", B"00110101", B"00100110", B"00010010",
 B"11011100", B"00100011", B"11100000", B"00101011", B"11001110",
 B"11101011", B"11101001", B"11010101", B"11011111", B"00111111",
 B"00011111", B"00001111", B"00100101", B"00100011", B"00100010",
 B"00101001", B"00101100", B"00110011", B"00011101", B"00000100",
 B"00101111", B"11100000", B"11011001", B"00010001", B"11001000",
 B"00010001", B"11101011", B"11001100", B"00001111", B"11100000",
 B"11011100", B"00100101", B"11011100", B"00100101", B"11010100",
 B"11000000", B"00110011", B"00101001", B"00101100", B"11100010",
 B"00111110", B"00111000", B"11101101", B"10101101", B"00100110",
 B"11110011", B"00010011", B"11011010", B"00001110", B"11001010",
 B"00110111", B"00010101", B"11101001", B"11100110", B"11011110",
 B"11110000", B"00010100", B"00010011", B"11100110", B"00100101",
 B"11101011", B"11101100", B"11001001", B"11011111", B"00100100",
 B"00011010", B"11011001", B"00010111", B"11100111", B"00101100",
 B"00001001", B"00101000", B"11101000", B"00110100", B"11011110",
 B"00010010", B"11110110", B"00011110", B"00101010", B"11000011",
 B"00000111", B"00101001", B"11001100", B"11011100", B"00101000",
 B"11101000", B"00110000", B"11011101", B"11100011", B"11000000",
 B"00101010", B"00100001", B"11110000", B"00110100", B"00110110",
 B"11011011", B"11110110", B"00100100", B"00011001", B"11001111",
 B"11001011", B"11000011", B"11100000", B"00001001", B"00000000",
 B"00011101", B"11011111", B"11101001", B"00111010", B"00100101",
 B"11001101", B"00110100", B"11011111", B"11001011", B"11111111",
 B"00110000", B"00101000", B"10111111", B"00011100", B"11100001",
 B"11101000", B"10111100", B"00011101", B"01000100", B"11100010",
 B"11001111", B"11111001", B"00100000", B"00010110", B"00100111",
 B"00101010", B"11100000", B"11011011", B"11101110", B"11110101",
 B"00010100", B"00010111", B"00011101", B"00011101", B"11001001",
 B"11011110", B"11101011", B"00111010", B"00001001", B"11110101",
 B"11100111", B"11011111", B"11011110", B"11001100", B"00101001",
 B"11101110", B"00101001", B"00000010", B"11101000", B"11100111",
 B"00110000", B"00010000", B"00100000", B"00010111", B"00110111",
 B"00100111", B"00101111", B"00000111", B"00100011", B"00010000",
 B"00101010", B"11101110", B"11100100", B"11101001", B"11010010",
 B"00011000", B"11010101", B"00001010", B"11011100", B"11100100",
 B"11010011", B"11111010", B"00000111", B"11111011", B"00101011",
 B"00010101", B"11111011", B"00000100", B"00110010", B"00100111",
 B"11010101", B"00010000", B"11010100", B"00110000", B"00101111",
 B"00111110", B"11100000", B"00010001", B"00011011", B"11010010",
 B"11111010", B"00010010", B"00010101", B"11101001", B"00000101",
 B"00011000", B"11101000", B"00011100", B"00010001", B"11000100",
 B"11101010", B"11011011", B"00101101", B"00011101", B"00010111",
 B"00011000", B"11011000", B"11001000", B"11010011", B"00011010",
 B"00011011", B"11100000", B"11100101", B"11101110", B"11111100",
 B"10111111", B"00010101", B"11101100", B"11001010", B"11001111",
 B"11100111", B"00100110", B"11100011", B"00011000", B"11101000",
 B"00101010", B"00010101", B"11010011", B"11101001", B"11110011",
 B"11101001", B"10111111", B"00100010", B"11101001", B"00011100",
 B"11001110", B"11011101", B"11101000", B"00100110", B"00001011",
 B"00110111", B"00001000", B"00011001", B"00101001", B"00100110",
 B"00110101", B"00101100", B"00011000", B"11110100", B"11010100",
 B"11011000", B"00010101", B"00100000", B"11011001", B"00011000",
 B"11001001", B"11010000", B"01000010", B"01000000", B"00011000",
 B"11010110", B"00100001", B"11100000", B"00010001", B"11001010",
 B"00010010", B"11011011", B"11010010", B"11101010", B"00011000",
 B"00010101", B"11111010", B"00100110", B"11010000", B"11110000",
 B"11011011", B"11011100", B"00100010", B"11011000", B"01000100",
 B"00011001", B"11011110", B"00011100", B"11011011", B"11100111",
 B"11100110", B"00010010", B"00001111", B"11011110", B"00100011",
 B"00011000", B"11001110", B"00000101", B"11100011", B"11001011",
 B"00000011", B"00011011", B"10110110", B"00100111", B"11110101",
 B"11100010", B"11000100", B"00010010", B"00101110", B"11111100",
 B"00000111", B"00011000", B"00001011", B"00100110", B"00101000",
 B"01000000", B"00110101", B"11101101", B"11100100", B"00010011",
 B"00110000", B"00011100", B"00101001", B"11011110", B"11010001",
 B"00101000", B"11110011", B"11010110", B"11100001", B"11101001",
 B"00010111", B"11011110", B"00111011", B"11101011", B"00010001",
 B"00101010", B"11100110", B"11111010", B"11011110", B"11101100",
 B"11001100", B"11100000", B"11101001", B"11100001", B"00101110",
 B"01000100", B"11001110", B"00011010", B"11101100", B"11011100",
 B"00011110", B"00011110", B"11101011", B"11110100", B"11100110",
 B"11110010", B"11110011", B"11110001", B"00001111", B"11101100",
 B"11011110", B"11010111", B"00111100", B"01000011", B"11001111",
 B"11011110", B"00110101", B"10111000", B"00001011", B"11011100",
 B"11011101", B"00101001", B"00011100", B"00000010", B"00000100",
 B"11110100", B"11001000", B"00110011", B"00010100", B"11100010",
 B"11010011", B"11001111", B"11011011", B"11111010", B"11011011",
 B"00001100", B"11110100", B"11000011", B"00100000", B"11110111",
 B"11101111", B"00100101", B"11100000", B"00100100", B"11010010",
 B"11101110", B"00111001", B"00111001", B"11001101", B"00110000",
 B"11101110", B"11110111", B"11010110", B"00001100", B"00100011",
 B"00000101", B"11000010", B"00011110", B"00000001", B"11001011",
 B"11111010", B"00011110", B"00011001", B"11010110", B"11011110",
 B"11101010", B"00110111", B"00010111", B"11011010", B"00011011",
 B"11010111", B"11001001", B"00110100", B"11011010", B"11110100",
 B"11100100", B"00010011", B"00110000", B"11011001", B"10111000",
 B"00001011", B"11101010", B"11101011", B"11100110", B"00011110",
 B"00011000", B"11100011", B"11101101", B"11101000", B"00011010",
 B"11011110", B"00101101", B"11011011", B"11101100", B"00000000",
 B"00100000", B"11100010", B"11101010", B"11010100", B"11011000",
 B"11111110", B"11001111", B"00101010", B"00100010", B"11011011",
 B"00010001", B"11010110", B"11001110", B"00000010", B"00011110",
 B"00100110", B"11101001", B"00111010", B"11110000", B"00111100",
 B"11010100", B"11011110", B"00011001", B"00110011", B"11110101",
 B"11101111", B"00100010", B"10111011", B"00001101", B"11011110",
 B"11110001", B"00011101", B"11000000", B"10111001", B"00110010",
 B"11011111", B"00110000", B"11001000", B"11011111", B"00000110",
 B"11011011", B"00100111", B"00010010", B"00011110", B"11010111",
 B"01001010", B"11101110", B"00101001", B"10111000", B"11010010",
 B"00011101", B"11110111", B"00110100", B"11100100", B"11010010",
 B"00011101", B"00011100", B"00101111", B"00001111", B"11010000",
 B"00111000", B"11011000", B"00100000", B"11100110", B"11001100",
 B"11010010", B"11001110", B"00110000", B"00101000", B"11100101",
 B"00101101", B"11110001", B"00101110", B"11010010", B"00011011",
 B"11100000", B"11010000", B"11010110", B"01000010", B"00110101",
 B"00011111", B"11100000", B"00110110", B"01001000", B"11110100",
 B"00010111", B"00100011", B"11100000", B"00011111", B"00011010",
 B"00000111", B"11100110", B"00100001", B"11101000", B"00010110",
 B"11011111", B"00011000", B"00100100", B"11100001", B"00100110",
 B"00011101", B"11010101", B"11110101", B"00101100", B"11101001",
 B"00000101", B"11011000", B"11100101", B"11100110", B"00100000",
 B"00000110", B"11110001", B"00000000", B"00100000", B"00110110",
 B"11011001", B"11010110", B"11100000", B"11011101", B"11010100",
 B"11001100", B"00100101", B"00110001", B"11100001", B"11101110",
 B"11010100", B"11011001", B"11101100", B"11100011", B"11100001",
 B"11010010", B"00100001", B"00010010", B"11110110", B"00011000",
 B"11011101", B"11010000", B"11011101", B"00001011", B"11011000",
 B"00011011", B"11100101", B"11010011", B"00100000", B"00100101",
 B"11110010", B"00001000", B"11100111", B"11100000", B"11010101",
 B"00010101", B"00011000", B"11111000", B"11011100", B"11110111",
 B"00101011", B"11001011", B"11101101", B"11011001", B"11001110",
 B"00101111", B"00101001", B"00001110", B"11100010", B"00011110",
 B"11011110", B"00000100", B"11100000", B"11011100", B"11100011",
 B"00001000", B"11010101", B"00010001", B"11011111", B"11010000",
 B"00010111", B"00011010", B"00110001", B"11101000", B"11011110",
 B"00001010", B"00000010", B"11101010", B"00000010", B"00010101",
 B"11001011", B"00000000", B"10111100", B"11011010", B"00111110",
 B"11101110", B"00001111", B"00010111", B"11100100", B"11001101",
 B"00110101", B"11011110", B"11010111", B"11010110", B"11110101",
 B"00101100", B"00110101", B"00011110", B"11101100", B"00100111",
 B"11111001", B"00011100", B"11010110", B"00010101", B"00010100",
 B"11010000", B"11101101", B"00011101", B"00000101", B"11100111",
 B"11100011", B"11011001", B"11110010", B"11011010", B"11101000",
 B"00011010", B"00101011", B"00000010", B"00000110", B"11111110",
 B"11011110", B"00010100", B"11101000", B"11010100", B"11100111",
 B"11111001", B"00110101", B"11011011", B"11011000", B"00100010",
 B"11001001", B"00011010", B"11101110", B"11010101", B"00111000",
 B"00000000", B"11100111", B"11101100", B"11010101", B"00011001",
 B"00001100", B"00100111", B"00010110", B"00001010", B"00101000",
 B"00101000", B"00100110", B"00010110", B"00101010", B"00101010",
 B"00101000", B"00000101", B"00011100", B"00110111", B"01000101",
 B"11100000", B"00100111", B"11010011", B"00010111", B"11100011",
 B"00010011", B"00110110", B"11010010", B"11110010", B"11100001",
 B"11110110", B"11110011", B"11100010", B"11011100", B"11101110",
 B"11110100", B"00011010", B"00101111", B"00100000", B"00001010",
 B"11011011", B"11111001", B"00101101", B"00111000", B"00011010",
 B"00100000", B"11101000", B"11100001", B"00101110", B"11111110",
 B"11001100", B"00011011", B"11011111", B"11000000", B"11011100",
 B"11101010", B"00010001", B"00101100", B"00010111", B"11010011",
 B"00101000", B"11110101", B"00100101", B"11011001", B"11011011",
 B"11111100", B"00110010", B"00011101", B"00100000", B"00011101",
 B"11011100", B"11101101", B"11010010", B"00101110", B"11100111",
 B"00010000", B"11001100", B"11110000", B"00100111", B"00011011",
 B"11100001", B"11000110", B"11011101", B"11110100", B"00101100",
 B"00001011", B"00101100", B"00011111", B"00011101", B"00100011",
 B"11011111", B"11100101", B"00010111", B"00101000", B"11011010",
 B"11101010", B"11000111", B"00100100", B"00110110", B"00001100",
 B"11010010", B"00101000", B"11100111", B"00100000", B"00001111",
 B"11010011", B"00010011", B"00101110", B"11000000", B"00111101",
 B"00000000", B"11110011", B"11011111", B"11010010", B"00100000",
 B"11110000", B"00100001", B"11100101", B"10111011", B"00010101",
 B"00111100", B"11010110", B"00011111", B"00010011", B"00000010",
 B"00010011", B"00110001", B"11101010", B"00011111", B"11110000",
 B"00101001", B"00101100", B"11010110", B"00101001", B"00010111",
 B"11111100", B"00000101", B"10111100", B"11100100", B"11100001",
 B"11011110", B"00001100", B"11010011", B"00011000", B"11010000",
 B"01001111", B"11101111", B"11111100", B"11010011", B"00100011",
 B"00101111", B"11101100", B"11011111", B"11100100", B"11011110",
 B"00100111", B"00110001", B"11110110", B"00110010", B"11101010",
 B"00000111", B"11101000", B"00001110", B"11010001", B"11100011",
 B"11110001", B"00010110", B"00001100", B"00110010", B"11010101",
 B"01000100", B"11110011", B"11011111", B"11110001", B"00101100",
 B"00101010", B"11000111", B"00110001", B"11001111", B"11011011",
 B"11100010", B"00011011", B"00110011", B"11110000", B"11111000",
 B"00011111", B"00011101", B"11010111", B"11011010", B"11011111",
 B"11001000", B"11111011", B"00011111", B"00010101", B"00001101",
 B"11100010", B"00101000", B"11101000", B"00000010", B"11101000",
 B"00001110", B"11100100", B"11001000", B"00000111", B"11001100",
 B"11110001", B"11010011", B"11100000", B"00101110", B"11010110",
 B"11011010", B"00110010", B"11111101", B"11010000", B"11101001",
 B"11100000", B"11101111", B"11010101", B"11101001", B"11111010",
 B"00001000", B"00110000", B"00010001", B"00001111", B"00000010",
 B"11010110", B"11011001", B"00101001", B"00100101", B"11101001",
 B"00100101", B"11001110", B"11100110", B"11100001", B"00100100",
 B"00001111", B"00010010", B"00011101", B"11011111", B"00010010",
 B"11111111", B"11101011", B"00100000", B"00101001", B"00111101",
 B"00100011", B"11011000", B"11111101", B"11001110", B"00011100",
 B"11001001", B"11011101", B"11100111", B"00011001", B"00001110",
 B"11000110", B"11100010", B"00100100", B"00011101", B"00001000",
 B"11110101", B"00110100", B"11011100", B"00101101", B"11100111",
 B"00110010", B"11101111", B"00010010", B"11110001", B"11110011",
 B"01000010", B"00011111", B"11000110", B"11001000", B"00101101",
 B"00111001", B"00010001", B"00100110", B"11100110", B"11011110",
 B"11001111", B"00001011", B"00111110", B"11101010", B"11010000",
 B"11011010", B"11010110", B"11111000", B"00100101", B"11000001",
 B"00100001", B"11011100", B"00000000", B"11110010", B"00001010",
 B"00101100", B"00101100", B"00010110", B"11111101", B"00101001",
 B"00010100", B"11111000", B"11010010", B"00011111", B"00110101",
 B"00101001", B"11111001", B"00100100", B"00100111", B"11011111",
 B"11111001", B"00101001", B"00101001", B"00110010", B"11100001",
 B"11100000", B"00100100", B"00110010", B"11011010", B"11100000",
 B"11011101", B"00100101", B"00101001", B"11100000", B"00010110",
 B"11101010", B"11001011", B"11010111", B"00011001", B"00001010",
 B"11101001", B"00100101", B"00011111", B"11010100", B"11001100",
 B"00110110", B"00011011", B"00010110", B"11110111", B"00110011",
 B"11110111", B"11110111", B"11100000", B"00011101", B"00000010",
 B"11010010", B"11000101", B"11111001", B"11100001", B"00001100",
 B"11011111", B"00110001", B"11001000", B"11100111", B"11010111",
 B"11101011", B"00000000", B"00001011", B"00011010", B"00101101",
 B"00010000", B"11011001", B"00011011", B"00100001", B"11101111",
 B"00101010", B"00101110", B"11100111", B"00101011", B"00011110",
 B"00000001", B"11101110", B"00011001", B"11000110", B"00111001",
 B"11100101", B"00111100", B"00011111", B"00001000", B"00010110",
 B"00010001", B"00010000", B"00100100", B"00111110", B"11100000",
 B"00100001", B"00010110", B"11111110", B"11100110", B"11010001",
 B"11101001", B"11011000", B"11010001", B"11101110", B"00110101",
 B"00101010", B"00101010", B"00011101", B"11100011", B"11100001",
 B"00000111", B"00100111", B"11011000", B"00011001", B"00001110",
 B"00000001", B"11011000", B"00101100", B"11100000", B"00001110",
 B"11100110", B"00011001", B"11110011", B"11101111", B"00011110",
 B"00010001", B"00100111", B"11100101", B"00101111", B"00100100",
 B"11100000", B"00011111", B"00110010", B"11110101", B"00011000",
 B"11101100", B"11101110", B"00101111", B"11101010", B"11010010",
 B"11010000", B"11011010", B"00100101", B"00011010", B"11101011",
 B"00011111", B"00111000", B"11011110", B"11111100", B"00100111",
 B"00011011", B"00111100", B"00101111", B"11100101", B"00101111",
 B"11011001", B"00100011", B"11101011", B"11011011", B"11111000",
 B"11101110", B"11010100", B"00100010", B"00001000", B"00001110",
 B"00010100", B"00100010", B"11100000", B"00100000", B"00100111",
 B"11010100", B"00100001", B"00110011", B"11100101", B"00110011",
 B"00010101", B"00100011", B"11001110", B"00100011", B"11001001",
 B"00110100", B"11001111", B"00011010", B"11011110", B"00110110",
 B"11100001", B"11110000", B"11010101", B"00100000", B"01000000",
 B"00111000", B"00110110", B"00011101", B"11001011", B"00100001",
 B"11010010", B"00100110", B"11010000", B"00100110", B"00011000",
 B"11001011", B"00011110", B"00001110", B"11100110", B"11010011",
 B"00001010", B"11110111", B"11110010", B"11101011", B"11100010",
 B"11110100", B"00101011", B"11010000", B"00001010", B"00110111",
 B"00100110", B"11010000", B"01001100", B"00001111", B"11100001",
 B"11011110", B"00101111", B"11010110", B"11000000", B"10110101",
 B"00010010", B"00101000", B"11001101", B"00010010", B"11110010",
 B"00100011", B"11100011", B"00011110", B"00011110", B"11001011",
 B"00110110", B"00101100", B"11101001", B"00101100", B"00100001",
 B"00100110", B"11001000", B"00100101", B"11011011", B"00110010",
 B"11101011", B"11100010", B"11011100", B"00111000", B"00101011",
 B"00111000", B"00100011", B"11100100", B"11100000", B"00001010",
 B"11011100", B"11100001", B"11111000", B"11101111", B"00011111",
 B"11010101", B"00111101", B"11111101", B"11101100", B"00100110",
 B"00001010", B"00100001", B"00101111", B"11111111", B"11100110",
 B"11010011", B"00100100", B"11011011", B"00011000", B"11101001",
 B"11011101", B"00011010", B"00100111", B"00101010", B"00100100",
 B"11100101", B"11011100", B"00011001", B"00010101", B"11100000",
 B"11100000", B"11100111", B"00001111", B"11011110", B"00110010",
 B"11011111", B"11100011", B"00101010", B"00010101", B"11011001",
 B"11100000", B"11100111", B"00101011", B"00100111", B"11101010",
 B"00011111", B"11011100", B"00101010", B"11011000", B"00111110",
 B"00110101", B"11010011", B"00110100", B"00100111", B"11111010",
 B"00100010", B"11101000", B"00111001", B"11000010", B"11010010",
 B"11000101", B"00100010", B"00101101", B"00001011", B"00110010",
 B"00010100", B"11010000", B"00100010", B"11011010", B"00010111",
 B"11001000", B"00110000", B"00101100", B"00110110", B"00110110",
 B"00010011", B"00101011", B"00101011", B"00110001", B"00011001",
 B"11010110", B"00010000", B"00100101", B"11100011", B"00101000",
 B"00000010", B"11011101", B"11001000", B"00100101", B"00010000",
 B"00101110", B"11101001", B"00101011", B"11100001", B"00010000",
 B"11011110", B"00110010", B"00101001", B"11100101", B"00000001",
 B"11100110", B"11111110", B"11101011", B"00011000", B"01000000",
 B"11101001", B"00100000", B"00100110", B"11010001", B"11100110",
 B"00101011", B"11111110", B"11011111", B"00101010", B"00011101",
 B"11011001", B"00000111", B"00011100", B"11101110", B"00111010",
 B"00011100", B"00111101", B"00001010", B"00111010", B"00100011",
 B"00101011", B"00011000", B"00010001", B"00001110", B"11010001",
 B"11011100", B"00110001", B"00011000", B"11110101", B"11110000",
 B"11011111", B"11010010", B"11011010", B"11001001", B"01000001",
 B"00100001", B"00111011", B"00110000", B"11011100", B"00101001",
 B"11011111", B"00011100", B"11110110", B"11101000", B"00100010",
 B"00110000", B"00010101", B"00011111", B"10111101", B"00011100",
 B"00110010", B"11011001", B"11101100", B"00010100", B"00110010",
 B"11101011", B"11010110", B"00100010", B"11100011", B"11001000",
 B"11110101", B"11010100", B"00011110", B"00001010", B"11101001",
 B"11011111", B"11000101", B"00011011", B"11001001", B"00100010",
 B"11110010", B"00000011", B"11000001", B"00110000", B"00111010",
 B"11100111", B"00111000", B"11011010", B"00011111", B"11100100",
 B"00111110", B"11100111", B"11100010", B"11001011", B"00101111",
 B"00011110", B"11100000", B"11110011", B"11011011", B"00001100",
 B"00101011", B"00100101", B"00100000", B"00010100", B"00101011",
 B"11010001", B"11100111", B"00011111", B"11010001", B"11100000",
 B"11010010", B"11001011", B"00011101", B"00011010", B"11101011",
 B"00101100", B"00011101", B"11101110", B"11111001", B"00110111",
 B"00100101", B"00001101", B"11010011", B"11100001", B"00101110",
 B"00101110", B"11011001", B"11101010", B"11010111", B"11100111",
 B"00010011", B"11100110", B"00101000", B"11001000", B"11001010",
 B"00100110", B"00101001", B"00100000", B"00100010", B"11101011",
 B"00100001", B"11000100", B"00111111", B"11011101", B"11100111",
 B"00000010", B"00001101", B"00110000", B"11100000", B"01000000",
 B"11101010", B"00101100", B"11101110", B"11010010", B"00100111",
 B"10111011", B"00100010", B"11101110", B"11011101", B"00100010",
 B"00110110", B"00001011", B"00100010", B"11001010", B"00010011",
 B"11000101", B"00010110", B"11011010", B"11110111", B"11100110",
 B"11100011", B"11010011", B"00011010", B"00100111", B"00001001",
 B"00011111", B"11101110", B"11010011", B"11101101", B"01000011",
 B"00011101", B"10111011", B"00011111", B"10111111", B"11111111",
 B"11101100", B"10111011", B"11010110", B"00101010", B"00011010",
 B"00010011", B"00101100", B"11011000", B"00011001", B"11110010",
 B"11011001", B"11101000", B"00110010", B"00110001", B"11001000",
 B"11101000", B"11111111", B"00000110", B"00010100", B"00000110",
 B"00011110", B"11010100", B"11111010", B"00100110", B"00100001",
 B"00100010", B"00000001", B"00011100", B"11011000", B"00111000",
 B"11101001", B"00011001", B"00110001", B"00001100", B"11101110",
 B"00010101", B"11010111", B"00011110", B"11101100", B"11011010",
 B"11010001", B"11100010", B"11110010", B"00010110", B"00001110",
 B"00101110", B"00100100", B"00010111", B"00010100", B"00011011",
 B"00011101", B"00010110", B"00100010", B"00101111", B"00100011",
 B"11011101", B"00010011", B"00011011", B"00110010", B"11100000",
 B"00101100", B"11001110", B"00001111", B"00100011", B"00101100",
 B"00100010", B"00100101", B"00100000", B"00110001", B"00100100",
 B"00010000", B"11011011", B"11010010", B"11010111", B"11011011",
 B"00101010", B"00010000", B"00011111", B"00101100", B"11011000",
 B"11100110", B"11010111", B"00011110", B"00011100", B"11111001",
 B"00100100", B"11010001", B"00010011", B"00100011", B"11100001",
 B"11010111", B"11111100", B"00011111", B"11010010", B"11011010",
 B"00101001", B"11011101", B"11010000", B"00100011", B"11101100",
 B"11011111", B"11100011", B"11100100", B"11101011", B"00001101",
 B"01000110", B"00101000", B"11011101", B"00100110", B"11001101",
 B"00101010", B"00100000", B"11100101", B"00011001", B"11011000",
 B"11010010", B"11100111", B"00011010", B"00010111", B"00011111",
 B"11111110", B"00001110", B"00101011", B"11101001", B"00110100",
 B"00111000", B"11100000", B"11100110", B"00100101", B"00001110",
 B"00001000", B"11011110", B"00011000", B"11010100", B"00100010",
 B"00100101", B"01000000", B"00010011", B"11100001", B"00100100",
 B"11100010", B"00001111", B"11010011", B"00100110", B"00011110",
 B"00001100", B"11111011", B"00100101", B"11010110", B"00001101",
 B"11101101", B"11100101", B"00011000", B"00100001", B"11011111",
 B"11100011", B"11000111", B"11010011", B"11001110", B"00010101",
 B"11010110", B"00100001", B"00110101", B"11101101", B"00001110",
 B"00100101", B"00000100", B"11000111", B"00011101", B"00011011",
 B"00111001", B"11000111", B"00100000", B"11100111", B"00100011",
 B"11101001", B"11101101", B"00110011", B"11001100", B"00001110",
 B"11000110", B"11111000", B"00001010", B"11111000", B"11011010",
 B"00100000", B"00100011", B"00010111", B"00111001", B"11001100",
 B"11110010", B"00011110", B"00011011", B"00101000", B"00101011",
 B"00010100", B"00010111", B"00101101", B"00100110", B"11010010",
 B"11100000", B"00010101", B"11000010", B"01000000", B"11001000",
 B"11000110", B"00100111", B"11000111", B"00001000", B"11010110",
 B"11111000", B"00101011", B"00110100", B"00101010", B"00000110",
 B"11000011", B"00010000", B"00000010", B"11000010", B"11010100",
 B"00011100", B"00111000", B"10111110", B"11101010", B"00011011",
 B"11110000", B"00000110", B"11110000", B"00111100", B"00101101",
 B"11101011", B"11101000", B"11101000", B"11110001", B"00001010",
 B"00101011", B"00001101", B"00011110", B"11011101", B"00000001",
 B"11100111", B"11110001", B"00011110", B"00100100", B"00011000",
 B"11010101", B"11100101", B"00011001", B"00000000", B"11011100",
 B"00100111", B"00110000", B"11100000", B"11100010", B"00010001",
 B"00111011", B"11101101", B"11010101", B"11100010", B"11010111",
 B"00010001", B"10110000", B"00010010", B"00010011", B"00110010",
 B"00101111", B"00010111", B"00011010", B"00010110", B"00011011",
 B"00011110", B"00101100", B"00100010", B"00101010", B"00110010",
 B"00101101", B"00110110", B"00001001", B"00110001", B"11011111",
 B"11010010", B"00100000", B"11010100", B"01000100", B"11100001",
 B"11010011", B"00110010", B"11010101", B"11011110", B"00110101",
 B"11100011", B"00010111", B"11010010", B"11100000", B"00010000",
 B"00001010", B"00100010", B"11110010", B"01000100", B"00001001",
 B"11011001", B"11110110", B"00100011", B"00011001", B"00101010",
 B"00001000", B"00100000", B"00011100", B"00010101", B"00101010",
 B"00100100", B"11010101", B"00011000", B"00011010", B"00110001",
 B"11110011", B"00001101", B"11001011", B"00110100", B"00111110",
 B"11100000", B"00111100", B"00110000", B"11011100", B"00011000",
 B"00101000", B"11110010", B"11010111", B"00111000", B"00100100",
 B"11010101", B"11001110", B"11011111", B"11000110", B"00000001",
 B"11101100", B"00001110", B"00010111", B"11011101", B"11110101",
 B"11100011", B"11101111", B"11001010", B"11110001", B"11011001",
 B"11100010", B"11110101", B"00100011", B"00011101", B"00011111",
 B"00101000", B"11100100", B"00001100", B"00011101", B"11011101",
 B"11100001", B"11000010", B"11101011", B"11100111", B"00011110",
 B"00100011", B"00000110", B"11000010", B"00011101", B"11100100",
 B"00011101", B"11011110", B"11011100", B"11101001", B"11011011",
 B"00101010", B"00011111", B"11000111", B"00101110", B"11111001",
 B"11000000", B"11010010", B"11100111", B"00000100", B"00111000",
 B"11011101", B"00010111", B"11010011", B"11011000", B"11000111",
 B"11010101", B"11100011", B"00100111", B"00010101", B"00011100",
 B"00101001", B"01000001", B"11100000", B"10110100", B"11011111",
 B"11101010", B"00110011", B"11011111", B"00011101", B"11000000",
 B"00110100", B"11110000", B"11101001", B"11100001", B"11010100",
 B"00011000", B"00110000", B"00110000", B"00101100", B"00001000",
 B"00101101", B"00100100", B"00101010", B"00000111", B"00100011",
 B"11110000", B"11001000", B"00100001", B"00110111", B"00000000",
 B"00101101", B"11101001", B"11100011", B"00010111", B"11100010",
 B"11100110", B"11100111", B"11100010", B"00100011", B"11101000",
 B"01001010", B"11110001", B"11011100", B"11001010", B"00011000",
 B"00101011", B"11110110", B"00100101", B"11010101", B"11100011",
 B"00011001", B"11001111", B"00010010", B"11010101", B"11110100",
 B"00101101", B"00101101", B"00100001", B"11011111", B"00100100",
 B"11110100", B"11100010", B"00100000", B"00011011", B"11101101",
 B"00110000", B"11010010", B"00001101", B"00110011", B"11000000",
 B"00011010", B"00110110", B"11100010", B"01000010", B"00110010",
 B"11101000", B"00100111", B"11101111", B"11110111", B"11001000",
 B"00010011", B"11100111", B"11001110", B"00110010", B"00000011",
 B"00011000", B"11011110", B"11001001", B"00100001", B"00100010",
 B"00011110", B"00010010", B"00100101", B"00011101", B"00111001",
 B"00001100", B"00010111", B"11010010", B"11000110", B"00010000",
 B"00100011", B"00101011", B"00000010", B"11010010", B"10111100",
 B"00100110", B"00001010", B"11101111", B"11010001", B"00010011",
 B"00101110", B"00001001", B"11101000", B"11011000", B"11100011",
 B"00100101", B"00001100", B"00010111", B"00111010", B"11110111",
 B"11010110", B"01000111", B"00100100", B"11001011", B"11111001",
 B"00100000", B"00100001", B"11010111", B"11101000", B"00001011",
 B"00011010", B"11000101", B"00001111", B"00001101", B"11100101",
 B"11011111", B"00110001", B"11101101", B"00010001", B"00100111",
 B"11101111", B"11011100", B"11100010", B"11010110", B"00000011",
 B"00010100", B"00100101", B"11100111", B"00011010", B"00011100",
 B"11110110", B"11010101", B"00011110", B"11110110", B"00100011",
 B"11111101", B"11100110", B"11101010", B"00101101", B"00100000",
 B"11100001", B"00010001", B"11001101", B"11011011", B"00011101",
 B"11101001", B"11000001", B"11101001", B"11000010", B"10110100",
 B"00011000", B"11011011", B"00011001", B"11100100", B"11100001",
 B"00010001", B"00110110", B"11110001", B"00100100", B"11011011",
 B"11110001", B"11010001", B"00101010", B"00011010", B"11010100",
 B"11100011", B"11011100", B"11110010", B"00001110", B"00010100",
 B"11101011", B"00010111", B"11011101", B"00011010", B"00010110",
 B"00100110", B"10111010", B"00010110", B"11010110", B"00110000",
 B"11101100", B"00110000", B"11110110", B"10110110", B"00110000",
 B"11010100", B"11100101", B"11100001", B"11010010", B"11011101",
 B"00001011", B"00100010", B"11001011", B"11110000", B"10111100",
 B"11011010", B"11011110", B"00011001", B"00001010", B"00100110",
 B"00010011", B"00100100", B"00000101", B"00100001", B"00010001",
 B"11000101", B"11100000", B"11110100", B"11011101", B"00000111",
 B"00010000", B"00100011", B"00001001", B"00101111", B"11011111",
 B"00110011", B"00110010", B"11011110", B"00010111", B"00110011",
 B"11100111", B"00100111", B"11100011", B"00011101", B"00011100",
 B"11110000", B"00111010", B"00100100", B"11101111", B"00011001",
 B"00010010", B"11100111", B"11110100", B"00001000", B"00101010",
 B"11010101", B"11100000", B"11010011", B"11001001", B"00010111",
 B"11110010", B"00100111", B"11100001", B"11100011", B"00000100",
 B"00011000", B"11011001", B"11100010", B"00001101", B"00010011",
 B"11110010", B"11101101", B"11011001", B"11010110", B"10110011",
 B"00101011", B"11001111", B"00101110", B"11110001", B"11100111",
 B"00011100", B"00010010", B"11100010", B"00100001", B"11110110",
 B"11110101", B"11101101", B"00100010", B"00101100", B"00011111",
 B"11111110", B"00110110", B"11011000", B"00100101", B"11010111",
 B"00111100", B"00000110", B"11100010", B"11100110", B"00011010",
 B"11111100", B"00100011", B"00001111", B"11011010", B"11011001",
 B"11100100", B"11110001", B"00010011", B"11100111", B"00010010",
 B"11011001", B"11111100", B"01010111", B"00011111", B"11100101",
 B"00100011", B"00111011", B"11100000", B"00010011", B"00101011",
 B"11101010", B"00010110", B"00011001", B"00001101", B"11010100",
 B"00101110", B"11101000", B"00100110", B"11000110", B"11001110",
 B"11011010", B"11100000", B"00011111", B"00011111", B"11101001",
 B"00010111", B"11101110", B"00010001", B"00010011", B"11011101",
 B"11101000", B"00010110", B"00100010", B"11010011", B"11001101",
 B"11101011", B"11010010", B"00101100", B"11100000", B"00011000",
 B"11100010", B"10111111", B"00101100", B"11100110", B"11010101",
 B"01001111", B"11000101", B"00101101", B"11010011", B"11100100",
 B"00010000", B"00000110", B"00011011", B"00100101", B"00110101",
 B"00100100", B"00010101", B"00010011", B"00111100", B"11011000",
 B"11101000", B"11000010", B"00010111", B"00101010", B"11010111",
 B"00001110", B"10111000", B"00100101", B"00110000", B"11001011",
 B"00010001", B"00010010", B"10110100", B"11011111", B"00010010",
 B"11101010", B"00011111", B"11111101", B"11010010", B"11100101",
 B"11001111", B"11000011", B"11100110", B"00100000", B"11101100",
 B"11110100", B"00011101", B"11100011", B"11100011", B"11100111",
 B"11100100", B"11011000", B"00011110", B"00100011", B"00001111",
 B"11101101", B"00010101", B"11011110", B"00100100", B"00011001",
 B"00010111", B"11111100", B"00010101", B"00100101", B"00011100",
 B"00100010", B"00001000", B"11101111", B"00011001", B"00010100",
 B"00101010", B"11110000", B"00001010", B"11110000", B"00011100",
 B"11000100", B"01010011", B"11010100", B"00110011", B"11110000",
 B"11011110", B"00010111", B"01000010", B"11011000", B"00100100",
 B"11101000", B"11011000", B"11011110", B"00111111", B"00011110",
 B"11010101", B"11010001", B"01001011", B"00011100", B"00101010",
 B"11001111", B"00111101", B"11010100", B"00011101", B"00010110",
 B"11101100", B"11100101", B"00011010", B"11100101", B"11011100",
 B"11100010", B"11000110", B"00011110", B"00100110", B"11101111",
 B"00101001", B"00100000", B"11110000", B"11011100", B"00010001",
 B"11001100", B"00111010", B"11100010", B"00000000", B"11011010",
 B"11011011", B"00100010", B"00010000", B"11011000", B"11100001",
 B"11111011", B"11011001", B"00110111", B"00100011", B"00100010",
 B"00101110", B"11001001", B"00011110", B"00100110", B"00100000",
 B"11010011", B"00101110", B"11100100", B"00010001", B"00011010",
 B"00111011", B"11100111", B"11000100", B"00101010", B"00101000",
 B"11100111", B"11011001", B"11101011", B"00101100", B"11011000",
 B"00100100", B"11101110", B"11110101", B"00111000", B"00001100",
 B"00010001", B"00001001", B"00101101", B"00100010", B"00110111",
 B"00111101", B"00110010", B"00010100", B"00101010", B"00101100",
 B"11011111", B"00100101", B"00101110", B"11110100", B"11010010",
 B"00101000", B"11101101", B"00011010", B"11101100", B"11101011",
 B"11101011", B"00101000", B"00111001", B"11010111", B"11001111",
 B"11101000", B"11011010", B"00111110", B"00000111", B"11011000",
 B"00010010", B"11011001", B"11011001", B"00011110", B"00100001",
 B"00010001", B"11010110", B"00001100", B"11000110", B"00111000",
 B"00011100", B"00000111", B"11001100", B"11001101", B"00110110",
 B"00101000", B"11100000", B"11000011", B"00100111", B"00000111",
 B"00011001", B"00110010", B"11101100", B"00101111", B"00100001",
 B"11111001", B"00011100", B"11100000", B"00101010", B"11011100",
 B"11100110", B"11010011", B"00100000", B"00100101", B"10111101",
 B"00100110", B"00010101", B"11100100", B"11100001", B"11011010",
 B"00000011", B"11010001", B"00100110", B"11010001", B"00011101",
 B"00100111", B"11100011", B"00110000", B"00001000", B"11101100",
 B"00001001", B"10111110", B"11011000", B"11100111", B"11010011",
 B"00101000", B"11001011", B"00111001", B"11101011", B"11011011",
 B"11001001", B"11111010", B"00101001", B"11010010", B"00000000",
 B"11000110", B"00011111", B"11010000", B"11011010", B"11001111",
 B"11011010", B"00100000", B"10111110", B"00001011", B"00010000",
 B"00100000", B"11010111", B"11101110", B"00001111", B"00010001",
 B"11100011", B"11010111", B"00010000", B"11110101", B"11101010",
 B"11101010", B"11010101", B"00001110", B"11110000", B"00110101",
 B"00010011", B"11101100", B"00011110", B"00011110", B"11111000",
 B"00011001", B"00101100", B"11011110", B"11010111", B"00000010",
 B"00101010", B"00110101", B"00010101", B"00000100", B"11101010",
 B"11100111", B"11011000", B"00011111", B"11100100", B"00100100",
 B"11001101", B"11111011", B"00011010", B"00011101", B"00000000",
 B"11010000", B"11101001", B"00110100", B"11001011", B"11000011",
 B"11011111", B"11100001", B"11010111", B"00110101", B"11101110",
 B"00000000", B"11101000", B"00011101", B"00011011", B"11001101",
 B"11001100", B"11100001", B"11010100", B"11101011", B"00110010",
 B"00100111", B"00011000", B"00101010", B"11100110", B"11110110",
 B"11101000", B"00011000", B"00011001", B"11100000", B"00011001",
 B"11010111", B"11101001", B"00101110", B"11001101", B"11011010",
 B"11100111", B"00101010", B"00101000", B"11011011", B"00001000",
 B"11001100", B"11110101", B"11010110", B"11101100", B"00010001",
 B"11100111", B"00001011", B"11111010", B"11110000", B"11111110",
 B"00100111", B"00100010", B"11100010", B"00010111", B"11011001",
 B"00100100", B"00100100", B"11011010", B"11100100", B"00010111",
 B"00101010", B"11100011", B"11110110", B"00101011", B"00010110",
 B"11100001", B"11100100", B"00001101", B"00110100", B"11101011",
 B"11110000", B"00010111", B"00010001", B"11010000", B"11011101",
 B"00100101", B"00010010", B"11010110", B"11110110", B"00100001",
 B"00100111", B"00010100", B"11011101", B"00101001", B"11011101",
 B"00110001", B"11010000", B"00111111", B"11111010", B"11100000",
 B"00011100", B"11101011", B"11010011", B"11110000", B"11100011",
 B"11010101", B"11111100", B"10111010", B"00011101", B"00101000",
 B"11000111", B"00100100", B"11110000", B"11100100", B"00001100",
 B"00101110", B"00110111", B"11000111", B"00000010", B"11010100",
 B"00011110", B"00100111", B"00010011", B"00010000", B"00101100",
 B"00011011", B"00011111", B"01001111", B"00010110", B"11010100",
 B"11010001", B"00101100", B"00001110", B"00011000", B"00011101",
 B"11101100", B"11010110", B"00010001", B"00101011", B"00011101",
 B"11100010", B"00011100", B"11101011", B"00011100", B"11010101",
 B"00100110", B"11011011", B"00011101", B"00101001", B"11001001",
 B"00001110", B"00011111", B"11001110", B"00001010", B"00011101",
 B"00001011", B"11100011", B"00100011", B"11010100", B"00001111",
 B"11011010", B"00010001", B"00101111", B"11001110", B"00011101",
 B"00011010", B"11000100", B"11011100", B"00010000", B"11011001",
 B"00110001", B"00101111", B"11101011", B"11110110", B"11101111",
 B"11011110", B"11100110", B"00011101", B"00011000", B"11011000",
 B"11110110", B"00110010", B"00001110", B"11110000", B"11011100",
 B"00010111", B"11011011", B"00111110", B"00100111", B"11100010",
 B"00001110", B"00011111", B"11011001", B"00001110", B"00111010",
 B"11011000", B"11110010", B"00000101", B"00011010", B"11011111",
 B"11100000", B"00010001", B"00000101", B"11001010", B"11010101",
 B"00000111", B"00100011", B"11001001", B"11101100", B"00101001",
 B"11110001", B"11100001", B"11011011", B"11010000", B"00101000",
 B"11100110", B"01001010", B"11011101", B"00011001", B"00110100",
 B"11101110", B"00010100", B"11001111", B"11101010", B"11011110",
 B"11100111", B"11110111", B"11011001", B"11011010", B"00010111",
 B"00101100", B"00010001", B"00101110", B"11110110", B"11011100",
 B"00101001", B"11010100", B"00001100", B"11010011", B"11101010",
 B"00110101", B"00111101", B"00110001", B"00001100", B"00101011",
 B"00011110", B"00000100", B"00100010", B"00101001", B"00011110",
 B"00011001", B"00011110", B"00001100", B"00100110", B"00011110",
 B"11111111", B"00100000", B"11101010", B"00011111", B"11101111",
 B"00001100", B"11001001", B"11101000", B"11110111", B"00100111",
 B"00101110", B"00010000", B"00100100", B"00011001", B"00010101",
 B"00010001", B"00011010", B"00110100", B"00011000", B"11110101",
 B"11011001", B"00111000", B"11101101", B"11101001", B"11010011",
 B"11010001", B"00000001", B"11110001", B"11011101", B"01001000",
 B"11010110", B"11100100", B"11100110", B"11100100", B"00011111",
 B"00111101", B"00101000", B"11011110", B"00011011", B"11011001",
 B"00011011", B"11010000", B"11010000", B"11111001", B"00101111",
 B"00100111", B"00010100", B"00010110", B"11011011", B"11100111",
 B"11010101", B"11011001", B"11100000", B"11011101", B"00001010",
 B"00011101", B"00010010", B"00101001", B"11101110", B"11110011",
 B"00010001", B"00101110", B"00010111", B"00010110", B"11100101",
 B"11101001", B"00110001", B"00010111", B"00010110", B"00011101",
 B"00011001", B"00100110", B"00100101", B"00001011", B"11000111",
 B"00001111", B"00100011", B"11100000", B"11110000", B"10111100",
 B"11100010", B"11101000", B"11011100", B"11100100", B"00100001",
 B"11101000", B"00101100", B"11000000", B"11001111", B"00100011",
 B"00100010", B"00010011", B"00110110", B"11110111", B"00011001",
 B"11011100", B"00100000", B"11100001", B"11001100", B"00100011",
 B"00111110", B"11010111", B"11111101", B"11101000", B"11100101",
 B"11100110", B"00010010", B"11011010", B"00101000", B"10111001",
 B"11100010", B"11100000", B"00100001", B"00010010", B"00100101",
 B"11011001", B"00111011", B"11011111", B"11011100", B"11100111",
 B"00011110", B"00101100", B"00010111", B"11100111", B"00010110",
 B"11110000", B"11011110", B"11011100", B"00100001", B"00011110",
 B"11011110", B"00011110", B"00100100", B"00010101", B"11010111",
 B"00101101", B"11101100", B"00101000", B"00101101", B"11011011",
 B"00010110", B"11011011", B"11011001", B"11101011", B"11111000",
 B"00100000", B"00100100", B"00011000", B"00110000", B"11011000",
 B"00011101", B"11000000", B"00100111", B"11011110", B"11001111",
 B"11101111", B"00101001", B"00111110", B"00010010", B"00110101",
 B"11111110", B"11100000", B"11011110", B"11001110", B"11110010",
 B"11011111", B"00111100", B"00010000", B"00001111", B"00001111",
 B"10111111", B"11000100", B"11110101", B"11101010", B"00010110",
 B"00110110", B"00100011", B"00100101", B"11010100", B"00100100",
 B"00001011", B"00010111", B"11010011", B"00100100", B"11111001",
 B"00101011", B"00000010", B"11011111", B"11110010", B"00100100",
 B"00110001", B"11011100", B"00011100", B"10111111", B"11011100",
 B"00101111", B"00011000", B"00100001", B"11110010", B"00010010",
 B"11101111", B"11101101", B"00100001", B"11100000", B"00011010",
 B"11100100", B"11011011", B"11010110", B"00001100", B"00000100",
 B"00101101", B"00100110", B"11011010", B"11001011", B"00001010",
 B"00001110", B"11100011", B"11001110", B"11011010", B"11011111",
 B"11100011", B"11101010", B"00010100", B"00101001", B"00010111",
 B"00001111", B"00001101", B"11010110", B"11011110", B"00011010",
 B"11101100", B"11000011", B"11010101", B"11101000", B"11011101",
 B"00100001", B"00101010", B"11110101", B"11011110", B"11011110",
 B"11100000", B"11001100", B"11010000", B"11111011", B"11110101",
 B"00101001", B"11011011", B"11100110", B"00111011", B"00001110",
 B"00001001", B"00011100", B"11010100", B"11010010", B"00100011",
 B"00110001", B"11110010", B"11011100", B"11011010", B"11011010",
 B"11111010", B"11011101", B"00011100", B"11000101", B"11010010",
 B"00010010", B"00000001", B"00100001", B"11010111", B"11001010",
 B"11001110", B"00010010", B"00010001", B"11101101", B"00010111",
 B"00100010", B"11100010", B"00001010", B"00110100", B"11110101",
 B"11111000", B"00100100", B"10111111", B"00000001", B"00100111",
 B"00011100", B"00010110", B"00101111", B"11110001", B"11011011",
 B"00100101", B"00011111", B"00011001", B"00110111", B"00100111",
 B"00100010", B"00011101", B"00100001", B"00101010", B"11001001",
 B"00100001", B"11100000", B"11100111", B"11010000", B"00010011",
 B"00010001", B"00011010", B"00011001", B"00100010", B"00100010",
 B"00100100", B"00011111", B"00110010", B"00100101", B"00011111",
 B"00100100", B"11101100", B"11101011", B"01000001", B"00011101",
 B"11101100", B"11011111", B"00001001", B"11010001", B"11011110",
 B"11111110", B"00110001", B"11001000", B"00010111", B"11011110",
 B"11110011", B"00101011", B"00001110", B"11100000", B"11010101",
 B"11110110", B"11011110", B"11000000", B"00010001", B"11100010",
 B"11011001", B"11011100", B"11110110", B"00100000", B"11100001",
 B"00001110", B"00111111", B"11110110", B"11000000", B"00001100",
 B"11100110", B"11110001", B"11011000", B"11101111", B"00101101",
 B"11100010", B"11111011", B"00100011", B"11100001", B"11011001",
 B"11010001", B"11110011", B"00100101", B"00111001", B"11100101",
 B"11100001", B"00011100", B"00110001", B"11111000", B"11101101",
 B"11001100", B"00001111", B"11000111", B"00101100", B"11110001",
 B"11100011", B"00011000", B"00001001", B"00100111", B"00010011",
 B"00010111", B"00001011", B"00011101", B"00100010", B"00011100",
 B"00010001", B"11011011", B"00101010", B"00100011", B"11111001",
 B"11001001", B"00011000", B"11010011", B"00101111", B"00001100",
 B"11100001", B"11110001", B"00000000", B"11101110", B"00101001",
 B"11011011", B"00101010", B"00001010", B"11110000", B"11011101",
 B"11101000", B"11011111", B"00100101", B"11101000", B"00100110",
 B"11010011", B"11011010", B"11101000", B"11101001", B"00100100",
 B"11000000", B"10110110", B"00011100", B"11110110", B"00010100",
 B"00101011", B"10111100", B"11111000", B"11100011", B"11001110",
 B"11101111", B"00001101", B"00010000", B"00100011", B"11110000",
 B"00011011", B"11101110", B"00100011", B"11010100", B"11011101",
 B"00110111", B"11100010", B"11110000", B"11011000", B"00010011",
 B"00110110", B"10110110", B"11011010", B"11000110", B"00111011",
 B"00011000", B"00100110", B"00010111", B"11001111", B"11011100",
 B"11101011", B"11000110", B"00100011", B"11000101", B"00101110",
 B"11010001", B"11111101", B"00011000", B"00010001", B"11010110",
 B"11011100", B"00101100", B"11111010", B"11010111", B"10111101",
 B"11100110", B"11101011", B"11100110", B"00011011", B"11011010",
 B"00111010", B"11001001", B"11011001", B"00100001", B"00100101",
 B"00001111", B"11001111", B"00011111", B"00100010", B"11101000",
 B"11100111", B"00011100", B"11010011", B"00011010", B"11011111",
 B"00100010", B"11100010", B"11010101", B"00010011", B"00001000",
 B"00010111", B"00111000", B"00100100", B"11110000", B"00100011",
 B"11101001", B"00010010", B"11011010", B"00011010", B"00000011",
 B"00001010", B"11100011", B"00101011", B"11100110", B"00010001",
 B"11100101", B"00000010", B"11011000", B"11101111", B"11011111",
 B"11100100", B"00011001", B"11011101", B"00100110", B"00001011",
 B"00111001", B"00111101", B"11100100", B"00011011", B"11101111",
 B"00011010", B"11110011", B"11001011", B"00010000", B"11100110",
 B"11010001", B"11100110", B"00000000", B"00010110", B"11011010",
 B"11001011", B"11101000", B"00100010", B"00111110", B"00100111",
 B"00011100", B"11011101", B"11100010", B"11011000", B"11101001",
 B"00011110", B"11010010", B"00100101", B"11111011", B"11011111",
 B"00111000", B"00011111", B"00011001", B"11010111", B"00011101",
 B"00011110", B"11010011", B"11011011", B"00111101", B"00110100",
 B"00010111", B"00000101", B"11100011", B"00101111", B"11011010",
 B"00100011", B"11011110", B"00010011", B"11100110", B"11010011",
 B"00001010", B"11011110", B"11101110", B"11011101", B"11101000",
 B"11101011", B"11101010", B"00110000", B"11111100", B"00100011",
 B"11101001", B"11101111", B"00010000", B"11100101", B"11110011",
 B"11010110", B"11111100", B"00100001", B"00011010", B"00010001",
 B"00101001", B"00100110", B"00000110", B"00010110", B"11110100",
 B"00011001", B"11010001", B"00010011", B"11110100", B"00100001",
 B"00101010", B"11001011", B"11010010", B"00100001", B"00100101",
 B"11001110", B"11101000", B"00000110", B"00011001", B"00111010",
 B"11110111", B"00110001", B"11101110", B"00100000", B"11010101",
 B"11110110", B"00101101", B"11111000", B"00101011", B"11011011",
 B"11010101", B"00100001", B"00100011", B"01001001", B"11101000",
 B"00100000", B"00001101", B"11010100", B"00011001", B"00101011",
 B"11111100", B"00011000", B"00101111", B"00101111", B"11010111",
 B"00000011", B"11111100", B"00100000", B"11110111", B"11110010",
 B"11010000", B"11011011", B"11100111", B"11110110", B"00001010",
 B"00010010", B"00101101", B"00111000", B"00001101", B"11101010",
 B"11101101", B"00011000", B"00100001", B"11101110", B"11001010",
 B"11010101", B"00100111", B"11010111", B"00101100", B"11001111",
 B"11101110", B"00011111", B"00100111", B"11010011", B"00100110",
 B"11100000", B"11101011", B"11100100", B"00010011", B"00110000",
 B"11011011", B"11001111", B"00110111", B"00001101", B"00010110",
 B"11100101", B"00110010", B"11110011", B"00011001", B"10111010",
 B"11100100", B"00100000", B"11100011", B"00011101", B"11010100",
 B"11100011", B"00110000", B"00011001", B"00000011", B"11110000",
 B"11111101", B"00110011", B"00100110", B"11100111", B"11100100",
 B"00111101", B"00010101", B"11011111", B"00101011", B"00011001",
 B"11100010", B"11010110", B"00101101", B"00011111", B"00100000",
 B"00101111", B"11100010", B"00100000", B"11001011", B"00010010",
 B"11100111", B"10111100", B"11010110", B"11010101", B"00010100",
 B"00011100", B"11010001", B"00110100", B"11011011", B"00100011",
 B"11010100", B"00011111", B"11011110", B"11010101", B"11111001",
 B"00011111", B"00100101", B"11100110", B"11000010", B"11110010",
 B"11010010", B"00011101", B"00011100", B"00011010", B"00110001",
 B"00000110", B"11100110", B"00011010", B"11111101", B"11011100",
 B"00000000", B"00101000", B"00100011", B"11100101", B"00010101",
 B"00100011", B"00101110", B"11011100", B"00110101", B"11100110",
 B"00100111", B"11011000", B"00100101", B"00101100", B"11101110",
 B"00000110", B"11101011", B"11010100", B"11011010", B"00010001",
 B"11100010", B"00100011", B"11100110", B"11100100", B"11011000",
 B"00100110", B"00001010", B"11101010", B"00011001", B"11100001",
 B"11011000", B"11001101", B"00010000", B"00110000", B"11101011",
 B"00110010", B"11001001", B"11011011", B"11100001", B"11101010",
 B"00100111", B"11010000", B"00100010", B"11010101", B"11110001",
 B"11011110", B"11011101", B"00011001", B"00111110", B"00010000",
 B"00101100", B"00001111", B"00110100", B"00010000", B"11101011",
 B"00100100", B"11011011", B"00000110", B"11010011", B"01001011",
 B"11101011", B"00100000", B"00001111", B"11101010", B"00101100",
 B"00100010", B"11111011", B"11011111", B"11100110", B"11100001",
 B"11000001", B"00110111", B"00011111", B"00101001", B"00101110",
 B"11101100", B"00110100", B"00100110", B"00010000", B"11101011",
 B"00001001", B"11011101", B"00011010", B"11110000", B"00011101",
 B"00011100", B"00000100", B"11100101", B"00011010", B"11101011",
 B"00010010", B"00010011", B"11011111", B"11010100", B"11001001",
 B"11011010", B"00100011", B"11010100", B"00101010", B"00111011",
 B"11001111", B"00000011", B"11010110", B"11001110", B"11010100",
 B"00010010", B"00101001", B"00101110", B"00000001", B"11101111",
 B"11011101", B"00101101", B"00001111", B"11110101", B"11101001",
 B"01000011", B"00010010", B"00101010", B"10110100", B"00011100",
 B"11011110", B"00100110", B"11001111", B"00001111", B"00001001",
 B"00011011", B"01001100", B"00101000", B"00011010", B"01001111",
 B"00010101", B"00001010", B"11100111", B"00110010", B"11000111",
 B"11101111", B"11010011", B"11111011", B"00011010", B"11101101",
 B"11011111", B"00101010", B"11001100", B"00011010", B"11100100",
 B"11011000", B"00011111", B"11100101", B"11011111", B"11011011",
 B"00001101", B"00001000", B"11111000", B"00110011", B"11001011",
 B"00110101", B"00011100", B"00101010", B"11100101", B"00001001",
 B"11100011", B"00000010", B"11001111", B"00011010", B"11011000",
 B"11101111", B"00010101", B"11100011", B"11110101", B"11010001",
 B"11010010", B"11010011", B"00001010", B"11010000", B"11000010",
 B"11000101", B"00001111", B"00001001", B"11110010", B"00011111",
 B"11011001", B"11100000", B"00110100", B"11100000", B"11100111",
 B"11010010", B"11010000", B"00101011", B"11101101", B"00001100",
 B"00011110", B"00100001", B"00110000", B"00100101", B"00011111",
 B"11011010", B"11100011", B"00000110", B"00110110", B"00100011",
 B"00011001", B"11110100", B"00000101", B"00001111", B"00011101",
 B"00010111", B"11000101", B"00101000", B"11000100", B"00100111",
 B"11001010", B"11110000", B"11011001", B"00010100", B"00011101",
 B"00000110", B"00110010", B"11011100", B"11010111", B"11001111",
 B"00000000", B"00010101", B"11110000", B"00110110", B"11100001",
 B"11000010", B"00000110", B"11100100", B"11100000", B"11100000",
 B"11110111", B"00111001", B"00010001", B"00011010", B"00110111",
 B"00101011", B"11101010", B"11100001", B"11001100", B"11011010",
 B"00100010", B"11011010", B"00110111", B"00100111", B"00101001",
 B"00010101", B"11011000", B"00010111", B"11011110", B"00011111",
 B"11100010", B"00101011", B"11100101", B"00100001", B"00011000",
 B"11011011", B"00100110", B"00000010", B"11011000", B"00110001",
 B"11101101", B"00111111", B"00110001", B"11100011", B"00111111",
 B"00100011", B"11001001", B"11101011", B"11011100", B"00100110",
 B"00000111", B"00010010", B"00010000", B"11101111", B"11100111",
 B"11101010", B"11101001", B"00011000", B"00100101", B"00100000",
 B"00100001", B"11010001", B"11011111", B"11111000", B"11100000",
 B"01000010", B"11011000", B"00100110", B"11100100", B"11100000",
 B"00010110", B"11110010", B"00110000", B"11000111", B"00100101",
 B"11101101", B"11111100", B"00100011", B"00101010", B"11100010",
 B"00101010", B"11110100", B"11010101", B"11101011", B"00110100",
 B"00011111", B"11101111", B"11101111", B"00010010", B"11110101",
 B"00011110", B"11111010", B"11001101", B"00110001", B"00000100",
 B"11010111", B"00010000", B"11011000", B"11011100", B"11101100",
 B"00010111", B"01001000", B"11110111", B"11000101", B"11000010",
 B"00101000", B"11100011", B"00000110", B"11010111", B"11110000",
 B"00011111", B"11110100", B"11110001", B"11111110", B"00010101",
 B"11110001", B"00011011", B"00010100", B"11111110", B"00000111",
 B"11100111", B"00001010", B"00110100", B"11101101", B"00101011",
 B"00101101", B"11101010", B"00010000", B"00110010", B"11110001",
 B"11000111", B"00001010", B"00001000", B"11110111", B"11100001",
 B"11010101", B"10111101", B"11111100", B"11101000", B"00011000",
 B"00101100", B"00100110", B"00001110", B"11011101", B"00011110",
 B"11100001", B"00001110", B"11010111", B"11000000", B"00101001",
 B"00100010", B"00100101", B"11100000", B"11110001", B"00100110",
 B"11101010", B"11100000", B"11100101", B"11101100", B"11111000",
 B"11111011", B"00010110", B"11101000", B"11011010", B"11100101",
 B"11010010", B"11011011", B"00000000", B"10011101", B"11010100",
 B"11011011", B"00011000", B"00110101", B"00110001", B"00011101",
 B"00110011", B"11011010", B"11101010", B"00011101", B"11011001",
 B"11001100", B"11101100", B"11011001", B"00010100", B"11010001",
 B"11101010", B"00001010", B"11010100", B"11100101", B"11101000",
 B"11011100", B"00011101", B"00010111", B"00110101", B"00100010",
 B"00001111", B"00011000", B"00100110", B"00001100", B"11111011",
 B"00010110", B"11100010", B"00101101", B"11111101", B"11010000",
 B"00010111", B"00011110", B"00110001", B"11010011", B"11011111",
 B"11011010", B"11100011", B"00100111", B"11011100", B"00101011",
 B"00000110", B"10110110", B"11110000", B"10111100", B"11111000",
 B"00011011", B"11011000", B"00101010", B"00010110", B"00100001",
 B"11001101", B"11010010", B"00011010", B"00011111", B"11101011",
 B"11110001", B"00010110", B"11011001", B"00011000", B"10111110",
 B"11101011", B"11011001", B"00100110", B"00010101", B"11101000",
 B"00100111", B"00011110", B"11011010", B"11100110", B"11001000",
 B"11001111", B"11110001", B"00111001", B"00100110", B"00100010",
 B"00100111", B"11110100", B"01001110", B"00011111", B"00011111",
 B"00100000", B"11100000", B"11100101", B"11001101", B"11000110",
 B"00011110", B"11000100", B"00101101", B"00101001", B"11000110",
 B"11001000", B"00111111", B"11111010", B"11100011", B"11111011",
 B"11011111", B"11101111", B"11101001", B"00100000", B"00001011",
 B"00100001", B"00100110", B"11101010", B"11111111", B"00100001",
 B"00110000", B"01000001", B"11110101", B"00110010", B"11011010",
 B"00001110", B"11001110", B"11100100", B"11001011", B"00101100",
 B"00011110", B"00011101", B"00101100", B"11101010", B"10111010",
 B"00000001", B"00010011", B"11111010", B"11111101", B"11100010",
 B"10111001", B"01000000", B"00110111", B"00110100", B"11111010",
 B"00100110", B"11101001", B"11100010", B"11010111", B"00010011",
 B"00110001", B"00100011", B"00110011", B"00100001", B"00010000",
 B"00011001", B"00100011", B"00010111", B"00100010", B"00010101",
 B"00111111", B"00000010", B"00111101", B"00010011", B"11100011",
 B"11100001", B"00010110", B"11011010", B"11001101", B"11010101",
 B"11010011", B"00001111", B"00111011", B"00100110", B"00111010",
 B"01000011", B"00011010", B"11100000", B"11110101", B"00011100",
 B"00011000", B"11100010", B"11101101", B"11011110", B"00100111",
 B"00010011", B"11011001", B"11100001", B"11101011", B"11001000",
 B"11010011", B"11011101", B"00111011", B"01000110", B"00100110",
 B"10111100", B"00100011", B"11011001", B"00101111", B"00101111",
 B"11000000", B"00001101", B"11101001", B"11011000", B"11101010",
 B"00100010", B"00100101", B"00010101", B"11110010", B"11101100",
 B"00000000", B"11010100", B"11111100", B"11001010", B"11010011",
 B"11100101", B"00010001", B"00111000", B"11010011", B"11010110",
 B"11101110", B"11010001", B"11101001", B"11010011", B"11110110",
 B"11011000", B"00010101", B"00001110", B"11100111", B"00110010",
 B"11010110", B"00100000", B"11110111", B"11101111", B"11100111",
 B"11100000", B"00011000", B"11100101", B"01001001", B"11101110",
 B"00010110", B"11011000", B"11010010", B"00001100", B"00001101",
 B"00100000", B"11011100", B"11011000", B"00110011", B"00001111",
 B"00011101", B"11011110", B"00110100", B"11010010", B"00010110",
 B"00010001", B"00000001", B"00001011", B"11011101", B"00001001",
 B"11010000", B"00011011", B"11101111", B"11000110", B"00011111",
 B"00101100", B"11100011", B"11101010", B"11010110", B"11000010",
 B"11101011", B"11110010", B"11100011", B"11011110", B"00110100",
 B"00100111", B"11110000", B"00101111", B"11110001", B"11100001",
 B"00100010", B"11011101", B"11100100", B"11011011", B"00010101",
 B"00100010", B"00000010", B"00101110", B"11001101", B"00101011",
 B"11011111", B"11110001", B"11011111", B"00111001", B"00101011",
 B"00101101", B"00111010", B"00101010", B"11011101", B"00100111",
 B"11100010", B"00011010", B"11010111", B"00000000", B"11011001",
 B"11100011", B"11111101", B"00110011", B"00100001", B"00001100",
 B"00110010", B"11010010", B"11011111", B"11100101", B"11010010",
 B"00101111", B"00100100", B"00100110", B"00101111", B"00011011",
 B"00110100", B"11011100", B"00011110", B"00001111", B"11001111",
 B"11111001", B"00110001", B"11011011", B"11011111", B"00100000",
 B"11000110", B"00100010", B"11010101", B"11111010", B"00001010",
 B"00101110", B"11111011", B"11001001", B"00011000", B"00011100",
 B"11111010", B"11010101", B"00101011", B"00010011", B"00001010",
 B"11111000", B"00011001", B"01001001", B"11101100", B"11101111",
 B"00011010", B"11111001", B"00101110", B"00010110", B"11011001",
 B"00011001", B"11110001", B"00110100", B"11110100", B"00000100",
 B"11011011", B"00101010", B"11110111", B"11011000", B"00010000",
 B"00010101", B"11101010", B"00011011", B"11011001", B"00100000",
 B"00001010", B"11010010", B"00111101", B"00100111", B"11101010",
 B"11010110", B"11101000", B"00100011", B"11101100", B"00101101",
 B"11100000", B"11011000", B"00110000", B"11101000", B"00010010",
 B"00100100", B"11011100", B"11010101", B"11000110", B"11111001",
 B"11100111", B"11010111", B"00110000", B"01000010", B"11000101",
 B"11100001", B"11001101", B"11100011", B"11110001", B"11110001",
 B"00001000", B"00010011", B"00100110", B"00111101", B"00011111",
 B"11011001", B"11010011", B"11110010", B"00100010", B"00101100",
 B"00010010", B"11100010", B"00010100", B"11011110", B"00011101",
 B"11100011", B"00010000", B"00100100", B"11001010", B"10111100",
 B"11000111", B"00000010", B"11010011", B"00100001", B"00000001",
 B"11100101", B"00101011", B"00100010", B"11000111", B"11011101",
 B"00011011", B"00011111", B"11011100", B"11110000", B"11110000",
 B"10111100", B"00100010", B"11101110", B"00110101", B"11100111",
 B"00101111", B"11010001", B"00001100", B"10111111", B"11001110",
 B"00011101", B"00101110", B"00011101", B"00010001", B"11011010",
 B"11100011", B"00100110", B"00101010", B"11110010", B"11001010",
 B"00011110", B"00011011", B"11000000", B"00001111", B"00011110",
 B"11011110", B"11111111", B"00011110", B"11101000", B"00010001",
 B"11111010", B"11100011", B"11010101", B"00100101", B"00100100",
 B"11100100", B"00110100", B"00010010", B"11011010", B"11001001",
 B"00011010", B"00011001", B"11101101", B"11111100", B"11111110",
 B"11100111", B"11001100", B"00000110", B"11010111", B"11010101",
 B"11101101", B"11110000", B"11100011", B"00001001", B"11100001",
 B"00010100", B"11100101", B"11010010", B"00101000", B"00011011",
 B"00100000", B"11010001", B"11101100", B"11100100", B"11110011",
 B"00101001", B"11010000", B"00101001", B"00010100", B"00011110",
 B"11011110", B"00000010", B"00011100", B"10111100", B"11100101",
 B"00101011", B"00100101", B"11110010", B"11101111", B"11010001",
 B"10111010", B"00010110", B"11100110", B"00010000", B"00010000",
 B"00101000", B"11011000", B"11011000", B"01000001", B"00100000",
 B"11010111", B"11100001", B"00100101", B"00111010", B"11101110",
 B"11011100", B"00100001", B"00000011", B"11100001", B"11101010",
 B"00000111", B"11100001", B"01000101", B"01000101", B"11100111",
 B"00011001", B"00011110", B"11101101", B"11001010", B"11010101",
 B"11001101", B"00101000", B"00100000", B"11101010", B"00111100",
 B"11000101", B"11110100", B"11001101", B"00000001", B"00100000",
 B"01000000", B"11111100", B"00001111", B"11100101", B"11101011",
 B"11110100", B"00101101", B"00001101", B"00100110", B"00011100",
 B"11111011", B"11010100", B"00100100", B"00110001", B"00101101",
 B"11010101", B"00101001", B"11101011", B"00110000", B"11101010",
 B"00010101", B"00001111", B"11100100", B"11100001", B"00111000",
 B"00100101", B"11010001", B"11101001", B"00010100", B"00100100",
 B"00010010", B"00001010", B"00100100", B"00101010", B"00001110",
 B"00100111", B"11001101", B"00101001", B"11001110", B"00010100",
 B"11110110", B"11010011", B"00111110", B"00010011", B"10110011",
 B"11100111", B"11011101", B"00101000", B"00011001", B"11010111",
 B"00011001", B"11011001", B"00100000", B"11111111", B"11100101",
 B"00100010", B"00010010", B"11000000", B"00010000", B"00011111",
 B"11011111", B"00100101", B"00110111", B"11100111", B"11011010",
 B"11000011", B"11110100", B"11100101", B"11001110", B"00100001",
 B"00011111", B"00101000", B"11110010", B"00100000", B"11001101",
 B"00000111", B"11010111", B"11101101", B"00101000", B"00100001",
 B"00011011", B"00110101", B"11100001", B"11111111", B"11001100",
 B"00001011", B"00101100", B"00101000", B"11011111", B"00011110",
 B"11000110", B"00010100", B"00101001", B"00100011", B"11100101",
 B"00101001", B"00011111", B"11111000", B"11011101", B"00001001",
 B"00100010", B"00101100", B"00011011", B"11010100", B"00011110",
 B"11100111", B"00011110", B"11011101", B"00000000", B"11010011",
 B"11000011", B"00100001", B"11000100", B"11101110", B"11101001",
 B"11011000", B"00101000", B"11010101", B"00101000", B"00011101",
 B"11011100", B"01000000", B"00001101", B"11011110", B"11010101",
 B"00100000", B"11101111", B"11011000", B"11010100", B"00110100",
 B"00010111", B"11101100", B"11110110", B"00100011", B"00100100",
 B"00101011", B"11001101", B"00100001", B"11101011", B"00010011",
 B"11001111", B"11101000", B"11000100", B"11100001", B"00101010",
 B"00101011", B"00010110", B"00011110", B"11010100", B"00100000",
 B"00100110", B"11111000", B"11011110", B"11100011", B"11110000",
 B"11110001", B"00010101", B"00100100", B"00110111", B"11110111",
 B"00011011", B"11001111", B"00100001", B"11110001", B"11001101",
 B"11110010", B"00001001", B"11000001", B"00100111", B"11010111",
 B"11010011", B"00011110", B"00101111", B"00100111", B"00010000",
 B"11101100", B"00111110", B"11100111", B"00010101", B"00000100",
 B"00010000", B"00111001", B"00110100", B"00101000", B"01000011",
 B"00110101", B"00100011", B"00011110", B"00100011", B"11101110",
 B"00010110", B"11100011", B"11101000", B"11100100", B"00001000",
 B"00001011", B"00011001", B"11010101", B"11100000", B"11100100",
 B"11011011", B"00011100", B"11100100", B"00010001", B"11100111",
 B"00010111", B"00101011", B"00000111", B"11101110", B"11010010",
 B"11001101", B"11100111", B"11010101", B"00110001", B"11110000",
 B"11100111", B"11100111", B"00110011", B"00111111", B"11001111",
 B"11000101", B"00001111", B"00011011", B"00101101", B"11101110",
 B"00011110", B"11010001", B"00110010", B"00011011", B"11101000",
 B"11010101", B"11011100", B"11100111", B"00110000", B"11010010",
 B"00001111", B"11100110", B"00010010", B"00011010", B"11010100",
 B"11010111", B"11001010", B"11001011", B"11011000", B"11011111",
 B"00101000", B"00010110", B"00101010", B"11101000", B"00011110",
 B"11001100", B"00100000", B"00011100", B"00001001", B"11101011",
 B"11100000", B"00010111", B"00100011", B"11010100", B"11011100",
 B"11010101", B"11100100", B"00001010", B"00011000", B"00011111",
 B"00010011", B"11011001", B"11101101", B"11010001", B"00110011",
 B"00010111", B"00100001", B"11001000", B"00011101", B"11111000",
 B"00101110", B"11100110", B"11010000", B"11100011", B"11001101",
 B"00011101", B"00101101", B"00101010", B"01001011", B"11110001",
 B"00001111", B"11100101", B"00110100", B"11010011", B"11011000",
 B"00000111", B"00100000", B"00100000", B"11100000", B"11101101",
 B"11111010", B"11111010", B"00101010", B"11101000", B"00100011",
 B"00111010", B"00111100", B"00001101", B"11110101", B"00011000",
 B"11011111", B"00001110", B"11011011", B"00010001", B"11101011",
 B"00010000", B"11101011", B"11110000", B"11101000", B"00000101",
 B"00110001", B"11101101", B"00100100", B"00010011", B"11010000",
 B"11100000", B"11100010", B"11011100", B"11100000", B"11111010",
 B"11001001", B"11100010", B"11011010", B"00101000", B"00000101",
 B"00101110", B"00011010", B"11010001", B"11111100", B"00100110",
 B"11011010", B"00101001", B"11100111", B"11100100", B"00100001",
 B"11101000", B"11111011", B"11100000", B"00110101", B"11011001",
 B"11010100", B"00101001", B"00110101", B"00011010", B"11011001",
 B"00001010", B"00100010", B"00000100", B"00100100", B"00011100",
 B"11100010", B"00011111", B"00100100", B"11010110", B"00000101",
 B"00010111", B"11001110", B"11110001", B"00001001", B"00010011",
 B"11001110", B"00011100", B"11000111", B"11101100", B"11010100",
 B"00100111", B"00011111", B"11010110", B"00101001", B"11101010",
 B"00010001", B"11011101", B"11111001", B"00010010", B"00100001",
 B"11111010", B"00100011", B"11100111", B"11100000", B"00000010",
 B"00010110", B"01000111", B"11110010", B"00110111", B"11100000",
 B"00011010", B"00100111", B"11111100", B"00001001", B"00110011",
 B"11011111", B"11010100", B"11101111", B"00010110", B"00101101",
 B"11010011", B"00101000", B"11011001", B"00111000", B"00010010",
 B"11110011", B"11110001", B"00100101", B"11011111", B"11010001",
 B"11100001", B"11011011", B"11001011", B"00001101", B"00101001",
 B"11100100", B"11100001", B"11000101", B"11100010", B"11001101",
 B"11100100", B"10111110", B"00001110", B"00010001", B"00011001",
 B"00011011", B"11011001", B"11100000", B"11111000", B"00011110",
 B"00101010", B"00010010", B"10111100", B"00101100", B"11100111",
 B"00001101", B"10111111", B"11001010", B"00100000", B"11111011",
 B"11111000", B"00100100", B"11010111", B"11011010", B"00011110",
 B"00111111", B"11010101", B"11010110", B"00100101", B"00110111",
 B"11101100", B"10111011", B"11100011", B"00110100", B"00011010",
 B"11010001", B"11100011", B"11110010", B"11000111", B"11000011",
 B"01000011", B"00100111", B"11010011", B"11011101", B"00011100",
 B"00011000", B"11110111", B"11101010", B"11111010", B"11011001",
 B"00101100", B"11011100", B"00101101", B"11100100", B"11100101",
 B"00110000", B"11011111", B"11010001", B"00010001", B"00010110",
 B"00100010", B"00111001", B"11011100", B"11011000", B"00010101",
 B"00011101", B"00101110", B"00100101", B"00011000", B"00010111",
 B"00011000", B"00011110", B"10111001", B"00100011", B"11001001",
 B"00111111", B"11000110", B"11110111", B"00011001", B"00000110",
 B"11011011", B"00100010", B"00111000", B"00100101", B"11010111",
 B"00110000", B"11010001", B"00100001", B"11100000", B"00011110",
 B"00110010", B"11010111", B"11011101", B"11010101", B"11100001",
 B"11101001", B"00000010", B"11001011", B"11001111", B"00000111",
 B"11011110", B"00101001", B"11011110", B"00100001", B"11001101",
 B"00101001", B"00100101", B"11100001", B"11011011", B"11110001",
 B"10111101", B"11001011", B"11100010", B"11110101", B"00001110",
 B"00011100", B"00110101", B"00111100", B"11101110", B"11101011",
 B"00111000", B"00011010", B"00001011", B"00011110", B"00010010",
 B"00011001", B"00001011", B"00001010", B"00110110", B"11011001",
 B"00011100", B"11010111", B"11000100", B"11100011", B"00110000",
 B"00101111", B"00000011", B"11100000", B"00110011", B"11010110",
 B"11001101", B"11100110", B"00010010", B"00100110", B"00010001",
 B"00001010", B"11001001", B"00011000", B"00011111", B"11001100",
 B"11100001", B"00110011", B"11001110", B"00010101", B"11001110",
 B"11001001", B"11011110", B"00000110", B"01001101", B"11101100",
 B"00010010", B"11111001", B"00111000", B"11011000", B"11000000",
 B"11001010", B"00011001", B"00010110", B"11011001", B"11110100",
 B"00100001", B"00110100", B"00011010", B"00111001", B"11100100",
 B"11101001", B"00011110", B"11101100", B"00010010", B"11100001",
 B"11010001", B"11001000", B"00011011", B"00100111", B"11100010",
 B"00101011", B"00010010", B"11111010", B"11010110", B"11110101",
 B"11000111", B"11010010", B"11011101", B"00101110", B"11010000",
 B"00100011", B"11010100", B"11000111", B"00011011", B"00100000",
 B"11110010", B"00110001", B"00010111", B"00011001", B"11111010",
 B"00100010", B"11011000", B"00100110", B"11001110", B"11010010",
 B"00110100", B"00010101", B"00011101", B"00100110", B"11000010",
 B"11000111", B"11010111", B"00001110", B"00100111", B"01001111",
 B"11101001", B"00100000", B"11010110", B"00110010", B"11100011",
 B"11100100", B"00100011", B"11101011", B"00100111", B"11010010",
 B"11011000", B"00110001", B"11000100", B"11101110", B"00100011",
 B"11100001", B"11111011", B"00000000", B"11110100", B"01000000",
 B"00101101", B"00101010", B"00110111", B"11100001", B"00011111",
 B"11100110", B"00011101", B"11011011", B"00100010", B"10101111",
 B"11100101", B"00011000", B"11000011", B"11001010", B"11011111",
 B"11011110", B"00110101", B"11110010", B"11010010", B"00100010",
 B"11010010", B"11011001", B"11111101", B"11101100", B"00000010",
 B"00001001", B"11110010", B"11010111", B"11011001", B"00101100",
 B"00010110", B"11100010", B"11101110", B"00101111", B"11000100",
 B"00101011", B"11101010", B"11101011", B"00100100", B"00001110",
 B"00110010", B"00011111", B"11011101", B"00100100", B"00110101",
 B"10101111", B"11011110", B"00001101", B"11011100", B"11100011",
 B"00011111", B"00011110", B"00100100", B"01000010", B"11011001",
 B"11001100", B"00101100", B"11001000", B"00000000", B"11110110",
 B"11100011", B"00101001", B"11011111", B"00100011", B"00011001",
 B"00000101", B"00000100", B"00011001", B"00010100", B"11010111",
 B"11100000", B"00001010", B"00001001", B"11110000", B"11100010",
 B"00011111", B"11101100", B"11100000", B"11001110", B"11011101",
 B"00011101", B"00011010", B"00000100", B"11010111", B"00100001",
 B"11100010", B"00011111", B"11010001", B"00111110", B"00100010",
 B"11101010", B"00101000", B"00011001", B"11011001", B"11101101",
 B"00011111", B"11101100", B"11011001", B"11100010", B"11001001",
 B"00001011", B"00110000", B"00010111", B"00100101", B"00101101",
 B"11011101", B"11100110", B"00110110", B"11100110", B"11001111",
 B"11010001", B"10111011", B"00011110", B"11011010", B"00011111",
 B"11010011", B"11101001", B"11010010", B"00100010", B"00100010",
 B"11101010", B"11000011", B"11100101", B"11011010", B"00100111",
 B"00100100", B"00010100", B"00010111", B"00101111", B"00101001",
 B"11001110", B"11111001", B"00101000", B"00010101", B"11011110",
 B"11110000", B"11100011", B"11100001", B"11100101", B"11111110",
 B"00000001", B"11100110", B"00011101", B"11010001", B"00110101",
 B"00110110", B"00110100", B"00011011", B"00000111", B"00011011",
 B"00010011", B"00001000", B"10111001", B"00111000", B"11110010",
 B"00011001", B"00000000", B"11100001", B"00010000", B"00000100",
 B"00010100", B"11101110", B"11101000", B"00010101", B"11000001",
 B"11011011", B"11010110", B"11000110", B"11001110", B"11011010",
 B"00101110", B"11111011", B"00101110", B"11001100", B"11111111",
 B"00000110", B"00010001", B"00011111", B"11010110", B"00001010",
 B"00101101", B"00001111", B"11100001", B"11001100", B"11110100",
 B"00101000", B"11101111", B"00110110", B"11010101", B"11100010",
 B"00011100", B"00101000", B"00000010", B"11011001", B"11110000",
 B"11010100", B"11101100", B"00100101", B"11101100", B"00011100",
 B"00011000", B"00011111", B"00110110", B"00110011", B"00010101",
 B"00000111", B"00010010", B"00100100", B"00100100", B"11100001",
 B"11110010", B"00110101", B"11001000", B"11011011", B"11100001",
 B"11101111", B"00101111", B"00010100", B"11011011", B"00100000",
 B"00010110", B"11110101", B"11101110", B"00001110", B"00110100",
 B"00100110", B"00100000", B"11100011", B"00001011", B"11100101",
 B"00011110", B"11011110", B"00010101", B"11011100", B"00110111",
 B"00100100", B"11011110", B"00100101", B"00100110", B"11001111",
 B"11011011", B"00001000", B"11100100", B"11100100", B"11011100",
 B"00100001", B"00100110", B"11010101", B"00100011", B"00010110",
 B"11110001", B"11111010", B"00011100", B"00101100", B"00000101",
 B"10111100", B"00010100", B"11001111", B"11001101", B"11110000",
 B"11100101", B"00010110", B"11001100", B"00110010", B"00011101",
 B"11110111", B"00100110", B"00101001", B"11100100", B"00011010",
 B"00100010", B"11100001", B"11011110", B"00010100", B"10111000",
 B"00011101", B"11011000", B"11001101", B"00111110", B"00100110",
 B"00010110", B"11101010", B"11010000", B"11010101", B"11011101",
 B"00011010", B"11100110", B"00000111", B"10111101", B"11010111",
 B"11101000", B"00100101", B"00100011", B"11100100", B"00011111",
 B"11100011", B"11110011", B"11011110", B"00011111", B"00110011",
 B"00110111", B"00101101", B"11100001", B"11111011", B"11000101",
 B"11010010", B"11001110", B"00101111", B"00100100", B"11110111",
 B"00110010", B"11011100", B"11011111", B"00000001", B"00100111",
 B"11100000", B"00010100", B"11100001", B"11110010", B"00101010",
 B"00011101", B"00111011", B"11010100", B"11010111", B"00100011",
 B"00011101", B"11000000", B"11011011", B"00101110", B"11001000",
 B"11100000", B"11110110", B"11001100", B"00011110", B"11001010",
 B"00011101", B"00101000", B"00100010", B"11011111", B"01000000",
 B"00010001", B"11100011", B"11000101", B"00110101", B"01000111",
 B"00100011", B"00011100", B"00100110", B"00010000", B"00010111",
 B"00010101", B"01000110", B"10111011", B"11101001", B"11011110",
 B"11000100", B"00010101", B"00000001", B"00011100", B"00000110",
 B"00100011", B"00010110", B"11110011", B"00100101", B"00011111",
 B"11100010", B"00000111", B"00001110", B"11110101", B"11001111",
 B"00101101", B"00101001", B"00101000", B"00000100", B"11100010",
 B"11011010", B"00011000", B"11010111", B"11101110", B"00101110",
 B"11101101", B"11010100", B"11110101", B"11100011", B"01000111",
 B"00000110", B"11110001", B"00011011", B"00000110", B"11110010",
 B"11110110", B"11100111", B"00011000", B"00100101", B"00101001",
 B"00101101", B"00011101", B"00011101", B"00001011", B"00001101",
 B"00010110", B"00111000", B"00010011", B"00110011", B"00011011",
 B"00011110", B"00101101", B"00001111", B"11000010", B"00111000",
 B"11111111", B"00001110", B"11010001", B"11100011", B"00011100",
 B"00110001", B"10111100", B"11011000", B"00010100", B"11101010",
 B"00001001", B"11011000", B"11100100", B"00011011", B"00101101",
 B"11010010", B"00111000", B"00110010", B"00000101", B"00100100",
 B"00110100", B"11101010", B"00000001", B"11011010", B"11100101",
 B"11111011", B"11111011", B"00000111", B"11100111", B"00011110",
 B"00100001", B"00100101", B"00110010", B"11011100", B"00101110",
 B"11010111", B"00000011", B"11110000", B"11110011", B"00010111",
 B"11011110", B"00010111", B"11101001", B"11100110", B"00100110",
 B"00011101", B"00100101", B"00011111", B"00101110", B"00010100",
 B"00101101", B"00010110", B"00101011", B"00100110", B"00011011",
 B"00100110", B"11100100", B"11100101", B"00101001", B"00010110",
 B"11100111", B"11101111", B"11100000", B"00100010", B"10111101",
 B"11110010", B"11101010", B"00000011", B"00010101", B"11001111",
 B"11100100", B"00100000", B"11010011", B"00101011", B"11011111",
 B"11100111", B"00111101", B"00011101", B"11010100", B"11010000",
 B"00110111", B"00010100", B"00011010", B"00001100", B"11101111",
 B"11001101", B"11011111", B"00001010", B"00101100", B"00011001",
 B"11000111", B"00110000", B"11110110", B"00010111", B"00010000",
 B"00000011", B"00100110", B"11001111", B"11011011", B"11101000",
 B"00010001", B"00011111", B"11010010", B"11000100", B"11011011",
 B"00110010", B"00100000", B"11011001", B"00010010", B"11000101",
 B"11011101", B"11100011", B"00010100", B"11010000", B"00000000",
 B"11011000", B"11011110", B"00010110", B"11100011", B"00100001",
 B"00100010", B"11100001", B"11010101", B"11011001", B"11010001",
 B"11100010", B"11011000", B"11101101", B"11101101", B"00011111",
 B"00100101", B"11010101", B"00111100", B"11010100", B"11011011",
 B"11011011", B"11101111", B"11011011", B"00100011", B"11111111",
 B"00101110", B"00001111", B"11011100", B"11101110", B"11001110",
 B"00100111", B"00100101", B"11010111", B"00110010", B"11000111",
 B"00110101", B"11001000", B"11000110", B"11101110", B"11100100",
 B"00100110", B"11000100", B"00101001", B"11010001", B"11100000",
 B"00011101", B"11010100", B"00010111", B"11011111", B"11100010",
 B"01000001", B"11100011", B"00110000", B"11110111", B"00100010",
 B"11011100", B"11011010", B"00011110", B"00111001", B"11001001",
 B"00011011", B"00011101", B"11101101", B"11100000", B"11101100",
 B"11011110", B"11011000", B"11011011", B"00110111", B"11010111",
 B"00010110", B"00000011", B"11011110", B"00010111", B"00010111",
 B"11100110", B"11100111", B"11011110", B"11101011", B"00111010",
 B"00101010", B"00001100", B"11110100", B"00101000", B"11011001",
 B"11000001", B"11101110", B"11010010", B"00011101", B"11010000",
 B"00100111", B"00101001", B"11010011", B"11101111", B"00010101",
 B"11000110", B"11110101", B"11101010", B"11011011", B"11011101",
 B"00100001", B"00000000", B"00001100", B"11100111", B"00011000",
 B"11010000", B"00011111", B"11100111", B"00110010", B"11100110",
 B"00101010", B"11011110", B"00001001", B"00101100", B"00011111",
 B"00101111", B"11111111", B"00001111", B"11001000", B"11100111",
 B"11010110", B"00101100", B"00110110", B"11101010", B"11010111",
 B"11100111", B"00011100", B"00011001", B"11100110", B"00011111",
 B"11010000", B"11010010", B"00000000", B"11010110", B"00101000",
 B"11010100", B"11010111", B"00110111", B"00100000", B"00101010",
 B"00100100", B"00010011", B"00110110", B"00101011", B"00010110",
 B"00101010", B"00011110", B"00010101", B"11101010", B"11100100",
 B"11100010", B"11110000", B"00110011", B"11011011", B"00101011",
 B"00100110", B"11011011", B"00000110", B"00010101", B"11011000",
 B"11011110", B"11100111", B"11101000", B"11010100", B"11011010",
 B"11100001", B"11010001", B"00101011", B"00011111", B"00001100",
 B"00011111", B"11011110", B"00101101", B"00011010", B"00000110",
 B"11000100", B"01000000", B"11110011", B"00010110", B"11010001",
 B"00101100", B"00001011", B"11101000", B"11101001", B"11101110",
 B"11000101", B"11100000", B"00100001", B"11101001", B"11110110",
 B"00100000", B"11010101", B"11011000", B"11010001", B"11001001",
 B"00001101", B"11010011", B"00001100", B"11001101", B"11100110",
 B"11101010", B"11111111", B"00100011", B"00100001", B"00011000",
 B"11101101", B"00001101", B"00110110", B"11010001", B"11001100",
 B"00011000", B"11011100", B"00110011", B"10110111", B"11111110",
 B"11010000", B"00101101", B"00011011", B"11010111", B"11101101",
 B"11010110", B"11000011", B"11111011", B"00011000", B"00100100",
 B"00010011", B"00010110", B"00100000", B"00100100", B"00101110",
 B"00010101", B"00011000", B"00111000", B"00101001", B"00001011",
 B"11011001", B"10111011", B"00110100", B"00111110", B"11100110",
 B"00101100", B"11110100", B"11100101", B"00101001", B"11101010",
 B"00010010", B"11100010", B"11011001", B"11101111", B"00100111",
 B"00010001", B"00101100", B"11001000", B"00011110", B"11011010",
 B"11101111", B"11110011", B"00101001", B"00100000", B"11100011",
 B"11110001", B"00100010", B"10111001", B"00010100", B"11100101",
 B"11011001", B"11101110", B"00011100", B"11011000", B"11001011",
 B"11111001", B"00000011", B"00001111", B"11110111", B"11111111",
 B"00100010", B"11010101", B"11011000", B"11011110", B"11001111",
 B"00101011", B"11010010", B"00011100", B"00010101", B"11100001",
 B"00111100", B"11000010", B"11010011", B"11011111", B"00111001",
 B"00101101", B"00001111", B"00011010", B"11111010", B"11010100",
 B"00011100", B"00101000", B"11011010", B"11001010", B"00110011",
 B"11011000", B"00100001", B"11101000", B"11001100", B"11101001",
 B"00011000", B"00000000", B"00101010", B"00100010", B"11001001",
 B"11101100", B"00001100", B"00110011", B"11111000", B"11100111",
 B"00101110", B"00100000", B"11011101", B"11011001", B"00110000",
 B"00010111", B"11001100", B"11011110", B"11111011", B"00011110",
 B"00001111", B"00000000", B"11110110", B"00010001", B"11111110",
 B"00001110", B"11011110", B"11010100", B"00100010", B"11110001",
 B"11111110", B"11111100", B"11100010", B"00101100", B"11001011",
 B"00011010", B"11101100", B"00000111", B"11100111", B"00110010",
 B"00101101", B"11100101", B"11110110", B"00011101", B"00101111",
 B"00100010", B"11101010", B"11111011", B"11100001", B"00011011",
 B"00101010", B"11011110", B"11111010", B"11101011", B"11011100",
 B"00011111", B"11010101", B"00110010", B"11111000", B"00101100",
 B"11101010", B"00100001", B"00000010", B"11100010", B"00011110",
 B"00011001", B"11011000", B"11101000", B"00001110", B"00010110",
 B"00101110", B"00110000", B"11101000", B"11001100", B"11100111",
 B"10111101", B"11100001", B"00100110", B"00011101", B"11100101",
 B"01001010", B"11111100", B"00110000", B"11010111", B"00010011",
 B"00011000", B"11101100", B"11111110", B"00100101", B"11000111",
 B"00011101", B"00000100", B"11100110", B"11011111", B"00011100",
 B"00110000", B"11110000", B"11101010", B"11010101", B"11011011",
 B"11101100", B"00100100", B"00101100", B"11101110", B"00011000",
 B"11011010", B"11010010", B"00011101", B"00101111", B"11000111",
 B"11101001", B"11101001", B"00000000", B"11000111", B"11100010",
 B"00011111", B"11110100", B"11011101", B"11101111", B"00110101",
 B"00011111", B"11010100", B"00000110", B"11011101", B"00010100",
 B"01000100", B"11100111", B"00111000", B"00100001", B"11110101",
 B"11110001", B"00101100", B"11100010", B"00100101", B"11101000",
 B"11011000", B"00001000", B"00001110", B"11101000", B"00001001",
 B"11111000", B"00100111", B"11101101", B"11011111", B"00001110",
 B"00110101", B"00011011", B"11010110", B"00010100", B"11111011",
 B"11101110", B"11001110", B"00011111", B"00011111", B"11010010",
 B"00101001", B"11111000", B"11100110", B"11011001", B"00100101",
 B"00000010", B"11100011", B"00110011", B"11010011", B"00101100",
 B"11010010", B"11011011", B"11100010", B"00100000", B"00100011",
 B"11011111", B"00010001", B"11011011", B"11001111", B"11011101",
 B"00100100", B"00101100", B"00001000", B"00101110", B"11011001",
 B"00011011", B"00010010", B"11100010", B"00110011", B"00010001",
 B"11011001", B"00010010", B"11110100", B"11100111", B"00100001",
 B"11100010", B"11100000", B"11111011", B"11001000", B"00110000",
 B"11001001", B"11101000", B"00001000", B"10100110", B"11110111",
 B"11110100", B"11010110", B"11010011", B"00011101", B"00000011",
 B"00100101", B"11011111", B"00100111", B"11010010", B"00010101",
 B"00010001", B"00011011", B"11110101", B"00011111", B"11101111",
 B"11110001", B"11010000", B"00010001", B"11001100", B"11001100",
 B"11011010", B"11000000", B"00010101", B"00100100", B"00111000",
 B"00001111", B"00010000", B"00100101", B"11011110", B"00010100",
 B"00001101", B"11011011", B"11101011", B"11111001", B"11011001",
 B"11010001", B"11100100", B"11010110", B"00100001", B"00100110",
 B"00111010", B"00101100", B"11011001", B"00111100", B"11011101",
 B"11110101", B"11001110", B"00101100", B"00100010", B"11001000",
 B"11010001", B"00010111", B"00011111", B"00101010", B"11110011",
 B"00101000", B"11010110", B"00001101", B"00100010", B"00100010",
 B"00100011", B"00101010", B"00010101", B"00111000", B"00110001",
 B"00001101", B"00100010", B"11100010", B"00010001", B"00100000",
 B"11110000", B"00001100", B"00010010", B"11101101", B"00110000",
 B"11101000", B"11100110", B"00010101", B"11101111", B"11110110",
 B"11000011", B"11010011", B"00011110", B"00100111", B"00111100",
 B"11011001", B"00011011", B"11010011", B"00001010", B"11010010",
 B"00110101", B"00011011", B"11011011", B"00011101", B"00011010",
 B"11110100", B"11110110", B"00100011", B"00110110", B"00000100",
 B"00000101", B"11111100", B"11111010", B"11100100", B"00010110",
 B"11101010", B"00101000", B"11101100", B"11010000", B"00001101",
 B"11110000", B"11100111", B"11001000", B"11001110", B"00110011",
 B"11010101", B"00101000", B"00111101", B"11100110", B"00000110",
 B"00011001", B"11011101", B"11101101", B"11011101", B"11010101",
 B"11000100", B"00100110", B"00011011", B"00101111", B"00100000",
 B"00101000", B"11011100", B"11011011", B"00100011", B"11111101",
 B"11100000", B"11100011", B"11010011", B"00011010", B"00010010",
 B"00101110", B"11010100", B"00010001", B"11011100", B"00110111",
 B"11011100", B"00011110", B"00101000", B"11011110", B"00100001",
 B"00001110", B"11011001", B"11101001", B"00110110", B"11010010",
 B"01000011", B"00011010", B"11110000", B"11000101", B"11100100",
 B"11111000", B"11000101", B"00000101", B"00100010", B"11101001",
 B"11000100", B"00111001", B"00101001", B"11101100", B"11010100",
 B"00101100", B"00010111", B"11110111", B"11100011", B"00110011",
 B"01000011", B"11001110", B"11011010", B"00011100", B"11100101",
 B"00100010", B"00111011", B"11010100", B"01001011", B"00010110",
 B"11010010", B"00011010", B"11010000", B"11001001", B"10110010",
 B"00000000", B"00011111", B"11101001", B"00011010", B"00110100",
 B"11010111", B"00100010", B"00110001", B"11001011", B"01000110",
 B"01000101", B"11100101", B"11100001", B"11111010", B"11011111",
 B"11110000", B"00011101", B"00011010", B"00111110", B"00100111",
 B"00001011", B"11010111", B"00001110", B"00010100", B"11110110",
 B"00101001", B"00010110", B"11011101", B"00110111", B"11110110",
 B"00100011", B"11000100", B"11001010", B"11010000", B"11110100",
 B"00011101", B"00110011", B"11011111", B"00101101", B"00101101",
 B"11011001", B"00100001", B"00011110", B"00001000", B"00000110",
 B"00111000", B"00010000", B"00100101", B"11101110", B"00110110",
 B"11110001", B"00101010", B"00100010", B"00011001", B"11101111",
 B"11001101", B"00001001", B"00010110", B"11100111", B"11010111",
 B"11011000", B"00100001", B"00011000", B"00010000", B"11110100",
 B"11111100", B"11001110", B"00001110", B"00101100", B"00010100",
 B"11110011", B"11100001", B"00100010", B"00110011", B"11111000",
 B"11001101", B"00110100", B"11011010", B"11100111", B"00010111",
 B"11100010", B"11110101", B"11100001", B"11101101", B"11100001",
 B"01000000", B"00101001", B"11100111", B"11100110", B"11011110",
 B"11110111", B"11010100", B"00000101", B"11010101", B"00111111",
 B"10111101", B"11011100", B"10101111", B"00001010", B"00000110",
 B"11100100", B"11110001", B"00000010", B"11101110", B"11011101",
 B"11011000", B"11011101", B"11110000", B"00001010", B"00010101",
 B"00011011", B"00111001", B"00010001", B"00101110", B"11100100",
 B"11111111", B"11001011", B"00100001", B"11001101", B"11101101",
 B"11011011", B"00010100", B"00110011", B"11010110", B"00110010",
 B"00010000", B"11101101", B"00010101", B"00000101", B"11011000",
 B"11100001", B"00011110", B"00011000", B"00110011", B"00011110",
 B"00100100", B"00101010", B"00101111", B"00101000", B"00011001",
 B"00000111", B"00000100", B"11100110", B"00011011", B"00110101",
 B"11101011", B"11100000", B"00010100", B"00010011", B"00011011",
 B"11011001", B"00100111", B"00011011", B"11001100", B"11011111",
 B"00011001", B"11110000", B"11101000", B"11011010", B"00011010",
 B"00100111", B"11111001", B"00100000", B"11001011", B"00111101",
 B"11110110", B"00001100", B"00010000", B"11101000", B"01000000",
 B"00101110", B"10111111", B"00010001", B"00011111", B"11100011",
 B"00100111", B"00001001", B"11011101", B"11100100", B"00001011",
 B"00011001", B"11010001", B"00010101", B"00100100", B"11110010",
 B"00100110", B"00010011", B"11101110", B"00011110", B"11100000",
 B"10111111", B"00100010", B"11100110", B"11000111", B"11101010",
 B"11010000", B"11101100", B"00100001", B"00001110", B"11110011",
 B"11011101", B"11011101", B"11101100", B"11110001", B"11001001",
 B"11100100", B"00011001", B"11100110", B"00101100", B"11001010",
 B"11110110", B"00111001", B"11011110", B"00100000", B"11010011",
 B"00001100", B"11100011", B"11010001", B"00010111", B"00100111",
 B"11111000", B"11010011", B"10111101", B"11101101", B"00100010",
 B"00111010", B"00010000", B"00010001", B"11100110", B"11110001",
 B"00110001", B"11100001", B"00000111", B"11011100", B"11001110",
 B"00101101", B"00100011", B"11011111", B"11001001", B"00001110",
 B"11110011", B"11000111", B"11100001", B"11111011", B"00001100",
 B"11010001", B"00001010", B"00010100", B"10110100", B"00100000",
 B"00101001", B"11010111", B"00001000", B"11011110", B"11010110",
 B"11100110", B"11101101", B"00100110", B"11100010", B"00010111",
 B"00010000", B"11101101", B"11011110", B"11101000", B"11000101",
 B"00010101", B"11101101", B"00000111", B"11101010", B"00110000",
 B"00001001", B"00011111", B"11100001", B"00001101", B"11100000",
 B"00100101", B"00110010", B"11100001", B"11000010", B"11111001",
 B"11010011", B"00100110", B"11101110", B"00000110", B"11100110",
 B"00100111", B"00010001", B"00011001", B"11010101", B"00011100",
 B"11010011", B"00010100", B"00010001", B"00110011", B"11001111",
 B"00001111", B"00001011", B"11001100", B"11000100", B"00110111",
 B"00010000", B"11011011", B"11001000", B"00111111", B"11110011",
 B"11010001", B"11001111", B"11010110", B"11111100", B"00101111",
 B"00100010", B"00111011", B"11110000", B"00101011", B"11100010",
 B"00010100", B"11101110", B"00101110", B"00011100", B"11101100",
 B"11011101", B"11100010", B"11101111", B"11101001", B"00011110",
 B"00001110", B"11100111", B"11100011", B"00001111", B"00010000",
 B"11000101", B"11010001", B"11100010", B"11010011", B"00100111",
 B"00110001", B"00101000", B"00101101", B"11010001", B"11100011",
 B"00001010", B"00001111", B"11011111", B"00101000", B"00110101",
 B"11100010", B"11010010", B"00111110", B"11101100", B"00101010",
 B"11100111", B"00001111", B"00011010", B"11010011", B"11100000",
 B"01000011", B"11111101", B"11100100", B"11001111", B"11011010",
 B"00110110", B"00011011", B"00001000", B"00011111", B"00010101",
 B"00011000", B"11101111", B"11010110", B"00101010", B"00101000",
 B"11011011", B"11100001", B"00011010", B"00101001", B"00010001",
 B"00011100", B"00011011", B"00110100", B"11111011", B"00010010",
 B"11011010", B"11011111", B"11101011", B"11100010", B"00100010",
 B"00101111", B"00010000", B"00001101", B"11010000", B"11001101",
 B"00010010", B"00011011", B"00001001", B"00011111", B"10111111",
 B"11101100", B"00001111", B"00010101", B"00111001", B"11100110",
 B"00001100", B"11101011", B"00100100", B"11100000", B"11100010",
 B"00010011", B"00111101", B"00101000", B"11101111", B"00011010",
 B"11100110", B"11110110", B"00011001", B"11111011", B"00010001",
 B"11011010", B"00011100", B"11011000", B"00100011", B"11100100",
 B"11001011", B"00010110", B"00101101", B"00011010", B"11100010",
 B"00110001", B"11100101", B"00110001", B"00001111", B"11011110",
 B"11010111", B"00101100", B"11011011", B"11100011", B"11100110",
 B"00001100", B"11100000", B"00110010", B"11010011", B"00100001",
 B"11010100", B"11101011", B"00011011", B"00110100", B"00001011",
 B"11000011", B"11011000", B"11101110", B"00011011", B"00010100",
 B"00010111", B"00011111", B"00001011", B"11111001", B"00011000",
 B"00011100", B"11110000", B"00100001", B"00100010", B"11100011",
 B"00100100", B"11000001", B"11001100", B"11011001", B"11011010",
 B"00110001", B"11110000", B"00011011", B"00101100", B"00011010",
 B"11101001", B"00101111", B"00011000", B"11101001", B"11100110",
 B"00111101", B"00100010", B"11111000", B"11010010", B"11011010",
 B"11101111", B"00100100", B"11100011", B"00001011", B"11011011",
 B"01001110", B"00101100", B"11111000", B"11100000", B"11101100",
 B"11110111", B"11011000", B"00101011", B"10110110", B"00000110",
 B"00011001", B"11011101", B"01001000", B"00110111", B"10111011",
 B"00100001", B"00001000", B"00000001", B"11110001", B"00011000",
 B"11110011", B"00011010", B"11101101", B"11101110", B"00011100",
 B"00100000", B"00011101", B"11100011", B"00110001", B"11101000",
 B"01000111", B"00011110", B"11101000", B"00011001", B"00010110",
 B"11100100", B"00110011", B"00100111", B"11010110", B"11110001",
 B"11001011", B"11011010", B"00110001", B"01000100", B"11100000",
 B"00100110", B"11011001", B"00100001", B"00011111", B"11100001",
 B"00100101", B"00100111", B"11010111", B"10111011", B"00110100",
 B"00000001", B"11011110", B"11011001", B"00010110", B"00010110",
 B"11100100", B"00011010", B"11011011", B"00100101", B"11101110",
 B"11110010", B"00100010", B"11000111", B"11101111", B"11110111",
 B"11011000", B"11110110", B"00100000", B"00010010", B"00001101",
 B"11110110", B"00011010", B"11100011", B"00101000", B"00010010",
 B"11011100", B"11110001", B"00010000", B"11111110", B"11010101",
 B"11001101", B"11010001", B"00010111", B"11010111", B"00001000",
 B"11011111", B"11011001", B"00000100", B"11011100", B"00011000",
 B"00010010", B"11101000", B"11110010", B"00011001", B"11100100",
 B"11011001", B"11101001", B"11001111", B"00101101", B"00110000",
 B"00010101", B"11110011", B"00011011", B"11101001", B"00000110",
 B"11101101", B"00000111", B"11011101", B"11101001", B"00100111",
 B"11000110", B"11100010", B"11101110", B"10110011", B"00101010",
 B"00011110", B"00100100", B"11011000", B"00010001", B"11010101",
 B"00011001", B"11100100", B"11011100", B"11100010", B"00011111",
 B"11101010", B"00100110", B"11101110", B"11011100", B"00110000",
 B"11110011", B"00100000", B"00001010", B"00110011", B"11110110",
 B"00101111", B"11111010", B"00111010", B"11111100", B"11111100",
 B"11101011", B"11100101", B"00011101", B"00101100", B"11111110",
 B"00110110", B"11011010", B"00101111", B"00100101", B"11001011",
 B"11000000", B"11101010", B"11011100", B"11110101", B"00110111",
 B"00100000", B"11011000", B"11100101", B"00100010", B"00011010",
 B"11010101", B"11101111", B"00011100", B"00110100", B"11010011",
 B"11100110", B"00101100", B"00101000", B"11100111", B"11101010",
 B"11010100", B"00100111", B"11101011", B"11101001", B"11011100",
 B"00100011", B"00010111", B"11100100", B"11101001", B"11001100",
 B"11010011", B"11011000", B"00101111", B"00011100", B"00011000",
 B"00011000", B"11111101", B"11101100", B"00010100", B"00111000",
 B"00100000", B"00000101", B"11110001", B"11101011", B"11010110",
 B"00010110", B"00011000", B"11101011", B"11011101", B"11101010",
 B"11001111", B"11010010", B"11100000", B"10111101", B"00011000",
 B"11101111", B"00011010", B"11011110", B"11010011", B"00110100",
 B"11101010", B"11101100", B"11101001", B"11111101", B"00001001",
 B"00101101", B"00000101", B"00011101", B"00100001", B"00100001",
 B"11100100", B"00110101", B"00001001", B"11011011", B"11101111",
 B"00101111", B"11101000", B"11101101", B"00100001", B"11100011",
 B"00010111", B"11101000", B"11010001", B"00010110", B"00011110",
 B"00011000", B"11000010", B"00001011", B"00110101", B"10110101",
 B"11011000", B"00101100", B"11011100", B"00011110", B"11101000",
 B"00110000", B"11001110", B"00000010", B"01000011", B"00101110",
 B"00110010", B"11110000", B"00110011", B"00010010", B"11010100",
 B"00100101", B"00011011", B"11100000", B"11010100", B"00011001",
 B"00101000", B"00101011", B"11000101", B"00101010", B"11001001",
 B"00001010", B"00010101", B"00100001", B"00000111", B"00011111",
 B"00110111", B"00110110", B"00010110", B"00000110", B"00100011",
 B"00010010", B"00010000", B"00101001", B"00100011", B"00100001",
 B"00100001", B"00001100", B"11100010", B"11110011", B"00011100",
 B"00010000", B"00011000", B"00110000", B"11001101", B"11000101",
 B"11110001", B"00100111", B"11100101", B"10111011", B"10111101",
 B"00101000", B"00010101", B"11001101", B"00101011", B"11011011",
 B"00011010", B"00001111", B"10111101", B"00100000", B"00011001",
 B"11001101", B"00100011", B"00010000", B"11010111", B"11011001",
 B"00110010", B"00010110", B"11110101", B"11001100", B"00100010",
 B"11100011", B"00101000", B"00011001", B"11010111", B"00101000",
 B"00011010", B"11011000", B"11111010", B"11111001", B"00011011",
 B"11100001", B"11010110", B"11111110", B"11101111", B"11011010",
 B"11110100", B"00011011", B"00110111", B"11010010", B"11010101",
 B"11011010", B"11110100", B"11011010", B"00100010", B"00011111",
 B"11010101", B"11011111", B"00011010", B"00000101", B"11111110",
 B"10111001", B"11011000", B"00011111", B"00100100", B"11100101",
 B"11011110", B"11010101", B"11110100", B"11001011", B"00010001",
 B"11101010", B"11100100", B"00101111", B"11111001", B"11000110",
 B"11000100", B"11100111", B"11100000", B"11100010", B"11011110",
 B"11101010", B"00101010", B"00100000", B"00101001", B"00010111",
 B"11101100", B"00110100", B"11011100", B"11101110", B"11101011",
 B"00100001", B"00110000", B"11011111", B"00101000", B"00011101",
 B"00111000", B"11101011", B"00110011", B"11110110", B"00100001",
 B"11000010", B"11010100", B"00110111", B"11100100", B"11011101",
 B"11011000", B"00100000", B"00011001", B"11100010", B"00010001",
 B"00101101", B"00101110", B"00110000", B"00100010", B"00100111",
 B"00100010", B"00100110", B"00011001", B"11001101", B"11011000",
 B"00000111", B"11100110", B"11100000", B"11100011", B"11100111",
 B"00010110", B"11101011", B"00101100", B"10111101", B"11010100",
 B"11110111", B"00010011", B"00101001", B"00011011", B"11100001",
 B"11001010", B"11100100", B"11100111", B"00100101", B"11100011",
 B"00011011", B"00000111", B"11110011", B"00100101", B"11111001",
 B"11101011", B"11100001", B"00110011", B"00100111", B"11010110",
 B"11100101", B"00001010", B"11001001", B"00100011", B"11010111",
 B"11100000", B"00011011", B"00011001", B"00011101", B"11100000",
 B"11101101", B"00010100", B"00110110", B"11101011", B"11100001",
 B"00110011", B"11010101", B"11101001", B"00010001", B"11110110",
 B"11001110", B"11011101", B"11011010", B"11100101", B"11001101",
 B"00010110", B"00100111", B"00100101", B"00010100", B"11101000",
 B"11010111", B"11010011", B"11101111", B"00010101", B"11001111",
 B"11011010", B"11110001", B"11101010", B"00000001", B"11011110",
 B"11011001", B"11100011", B"00101001", B"00011011", B"11001100",
 B"00010010", B"11010001", B"11101010", B"11001101", B"11101111",
 B"11111000", B"00100101", B"00010111", B"00100011", B"00000111",
 B"11101101", B"11010111", B"00101001", B"11101010", B"00001101",
 B"11110110", B"11011011", B"00011001", B"00110000", B"11100001",
 B"11100100", B"00100110", B"11011101", B"11111010", B"11101101",
 B"11101010", B"11101010", B"00010000", B"11100110", B"00001100",
 B"11011011", B"11011000", B"01000000", B"00010110", B"00001111",
 B"11110100", B"00110000", B"11010011", B"11100111", B"11110010",
 B"00011111", B"00011101", B"11011011", B"00010011", B"00001100",
 B"00011111", B"11111010", B"00100100", B"11011111", B"00011001",
 B"11110100", B"00001000", B"11110110", B"00100010", B"11001101",
 B"11100001", B"00110110", B"00101000", B"00011011", B"00011100",
 B"00011001", B"00110000", B"00011101", B"00001001", B"00111010",
 B"00000011", B"11010111", B"00110010", B"11010001", B"11011111",
 B"11101010", B"00110100", B"00100110", B"11011010", B"11011001",
 B"11100100", B"00001100", B"00011100", B"00010111", B"00011110",
 B"11010010", B"11011100", B"11101010", B"00001000", B"00010101",
 B"00100110", B"11110100", B"00101100", B"11010100", B"00110010",
 B"11101000", B"11010010", B"11110001", B"11010101", B"00110111",
 B"00011100", B"00100101", B"00011010", B"00111011", B"11011010",
 B"00101100", B"11011001", B"11011010", B"11100011", B"00101010",
 B"00010001", B"00011111", B"11110000", B"11010010", B"11100100",
 B"11110101", B"00010111", B"11000100", B"00111001", B"11100101",
 B"00011000", B"11101011", B"11010011", B"11110110", B"00100101",
 B"00101000", B"11100000", B"00001001", B"11101001", B"00010100",
 B"11101111", B"11010011", B"11101111", B"00101000", B"00011111",
 B"10111111", B"11110011", B"00010011", B"11011101", B"00110011",
 B"11010010", B"11011110", B"00011101", B"11100010", B"11001101",
 B"11100001", B"00011000", B"00001111", B"11100011", B"00100101",
 B"11100110", B"01001101", B"11110100", B"00100111", B"11100011",
 B"11011001", B"11011110", B"00010101", B"00110010", B"11010110",
 B"00100101", B"00000110", B"00010111", B"11101100", B"00011000",
 B"11100001", B"00001101", B"00100010", B"00100111", B"11011111",
 B"11011100", B"00101001", B"00101101", B"00000000", B"11010101",
 B"11010010", B"11011011", B"00111100", B"11011011", B"00110110",
 B"11100001", B"11001110", B"00111011", B"11011111", B"00001100",
 B"11100001", B"00011111", B"00101110", B"11111000", B"00101101",
 B"11100101", B"00101110", B"11010111", B"10111100", B"00000101",
 B"11011111", B"11011111", B"11001011", B"11011001", B"11010000",
 B"11011111", B"00001011", B"00100001", B"00110010", B"00101010",
 B"11101000", B"11011000", B"11011110", B"11100011", B"11001100",
 B"00110100", B"00001000", B"11011110", B"00100011", B"11100010",
 B"00100001", B"00100010", B"00110000", B"00100001", B"00011001",
 B"00010100", B"00100000", B"00011101", B"11101101", B"00101000",
 B"11110100", B"11100110", B"11101000", B"00100100", B"00011001",
 B"11100000", B"11100011", B"00100101", B"11010001", B"11111100",
 B"11001101", B"00011101", B"00010110", B"11011010", B"00001011",
 B"00100010", B"00110001", B"00100101", B"00010101", B"11111010",
 B"00010100", B"00011110", B"00101001", B"00011100", B"00010011",
 B"11100001", B"00001111", B"11011111", B"00011111", B"11100101",
 B"00110111", B"00101100", B"11001011", B"11010111", B"00011111",
 B"00100101", B"11011001", B"11100101", B"11010011", B"11110011",
 B"00001110", B"11100110", B"00011010", B"11101110", B"11010001",
 B"00011010", B"00011110", B"00110111", B"11110101", B"11011100",
 B"00000111", B"00110001", B"11101001", B"00000101", B"11110011",
 B"11100101", B"11100011", B"11011111", B"00100000", B"00110010",
 B"00011110", B"00110000", B"11100000", B"00011101", B"00110111",
 B"00001111", B"11101001", B"00100010", B"11010110", B"00010110",
 B"11101101", B"11010010", B"00100011", B"11010110", B"00101011",
 B"11011000", B"11100011", B"00110101", B"11011011", B"00011100",
 B"00001101", B"11010000", B"11101001", B"11101000", B"11110001",
 B"11010011", B"11011101", B"11101100", B"11011110", B"00000001",
 B"00110101", B"11011101", B"00011110", B"11101011", B"11001010",
 B"11101001", B"00101110", B"00100011", B"00110010", B"00101010",
 B"11001010", B"11001100", B"00101110", B"11101111", B"00011101",
 B"00000111", B"11100110", B"00111010", B"00101000", B"11110001",
 B"00011001", B"11011100", B"11100100", B"11100011", B"11011001",
 B"00001100", B"11011001", B"00011010", B"00101011", B"00011011",
 B"11101000", B"00110001", B"00011010", B"11110000", B"11110110",
 B"00000111", B"00010111", B"00100010", B"11100100", B"00010100",
 B"00011001", B"11110011", B"11100110", B"00001110", B"11110000",
 B"00100100", B"00110101", B"11010110", B"11011100", B"11010110",
 B"11010011", B"11010101", B"00101101", B"11011110", B"11011011",
 B"11100000", B"11011101", B"00010100", B"11001100", B"00100010",
 B"11100000", B"11011111", B"00011010", B"11011010", B"01000111",
 B"11110001", B"11100101", B"00010110", B"00100110", B"11001000",
 B"00101100", B"11100100", B"11100001", B"11001110", B"11111101",
 B"00100110", B"00100100", B"11111110", B"00100110", B"00001110",
 B"11101000", B"00110101", B"00101110", B"11101010", B"00100011",
 B"00110100", B"11011000", B"00100010", B"00101101", B"11010011",
 B"11000111", B"00100011", B"11010111", B"00011001", B"00011100",
 B"00011100", B"11101100", B"00110000", B"11011010", B"11110110",
 B"11101101", B"00001101", B"00001100", B"00101000", B"00011110",
 B"00101001", B"00010101", B"00010101", B"11100010", B"00001100",
 B"00011110", B"11100001", B"11010110", B"11010011", B"11110111",
 B"11001100", B"11101010", B"00101111", B"11110010", B"11100010",
 B"11010101", B"00100000", B"00001000", B"11011001", B"00100010",
 B"11101011", B"11100001", B"00110100", B"11001000", B"11101001",
 B"11000011", B"11010001", B"11100110", B"11011110", B"11010010",
 B"00101010", B"00001111", B"11001011", B"00011101", B"11101101",
 B"00100001", B"11100101", B"00101011", B"00101100", B"11100110",
 B"00100100", B"00010110", B"11010110", B"00110110", B"00010011",
 B"11010101", B"11100101", B"00111001", B"00010111", B"11101000",
 B"00000001", B"11100110", B"11101101", B"00011100", B"00100110",
 B"00100110", B"00101101", B"11101000", B"11001010", B"00101000",
 B"00001111", B"00010001", B"11101010", B"00100111", B"11011011",
 B"00001000", B"11100101", B"00011001", B"11011100", B"11011110",
 B"11111010", B"11101111", B"00110001", B"11011010", B"11111111",
 B"00100110", B"00101100", B"00010101", B"01000011", B"00101011",
 B"01000010", B"00110100", B"00001011", B"11100010", B"00010011",
 B"01000100", B"11101000", B"11100011", B"11001000", B"11100011",
 B"11101101", B"11011010", B"11010001", B"00110000", B"11011100",
 B"00101111", B"11000111", B"11000001", B"00110000", B"11111111",
 B"00101000", B"00101000", B"00010000", B"01000101", B"00100001",
 B"00010010", B"00100000", B"11110111", B"11100011", B"11110010",
 B"11010011", B"00101100", B"00101000", B"00100011", B"00101110",
 B"00011001", B"00010111", B"11010100", B"11101111", B"00000110",
 B"00100101", B"11011001", B"11101001", B"11011001", B"00101000",
 B"00100101", B"00101101", B"11110101", B"00111010", B"11010101",
 B"11110100", B"11100011", B"00010101", B"11100001", B"11010100",
 B"11100011", B"00101101", B"00101111", B"11100011", B"00100001",
 B"00001101", B"00111010", B"11011110", B"00110110", B"11100000",
 B"00101001", B"11110101", B"00101010", B"11110101", B"00100011",
 B"11011100", B"11101110", B"11010010", B"00101001", B"00000000",
 B"00101001", B"00101010", B"00100000", B"11110011", B"11111011",
 B"11001010", B"00101011", B"11010110", B"11110011", B"11110110",
 B"11011001", B"01000001", B"00111001", B"11110010", B"00110100",
 B"10111000", B"11100110", B"11010111", B"00001110", B"00001111",
 B"00100001", B"00110101", B"11011001", B"11101111", B"00100101",
 B"10110111", B"00110100", B"11010001", B"11101100", B"11100000",
 B"00101110", B"00001100", B"11000101", B"11010111", B"11110011",
 B"00101011", B"00100101", B"11110110", B"00011100", B"11010100",
 B"00001111", B"00000000", B"11100111", B"00110011", B"11010011",
 B"11101110", B"11010001", B"11100110", B"00110100", B"00101000",
 B"11100000", B"11100010", B"00100001", B"00101000", B"11011110",
 B"00000100", B"00000010", B"11101011", B"00100000", B"00001100",
 B"11110010", B"00011000", B"00111110", B"11001110", B"00010011",
 B"11110010", B"00111100", B"11101000", B"11011100", B"11011101",
 B"00000001", B"00110101", B"00001110", B"11010111", B"11010110",
 B"11001110", B"11111101", B"00011010", B"00100000", B"00001110",
 B"00000101", B"11110101", B"11100101", B"00010100", B"11101100",
 B"11011111", B"00001100", B"11101001", B"00101001", B"11100100",
 B"00100100", B"11011010", B"11011110", B"11011101", B"00001001",
 B"00001000", B"00110000", B"00011111", B"11011000", B"10101101",
 B"00011110", B"00000111", B"11110011", B"11110110", B"11010101",
 B"00001001", B"11011100", B"11011011", B"11101110", B"00000001",
 B"00101000", B"11010001", B"00010110", B"11011110", B"00010111",
 B"00101011", B"11111101", B"00110100", B"00101001", B"11010010",
 B"11110010", B"11011100", B"11111100", B"00100111", B"00111001",
 B"11101001", B"00110001", B"11101010", B"00011000", B"00000001",
 B"11110001", B"00011111", B"11011000", B"11011110", B"11011010",
 B"11110011", B"11010000", B"11100111", B"00011101", B"00011110",
 B"00001110", B"00011000", B"11100110", B"11010101", B"11010000",
 B"00100111", B"11101011", B"00001111", B"10111001", B"11110101",
 B"00000010", B"00100001", B"00011010", B"11100010", B"11010101",
 B"11000011", B"11010111", B"00101101", B"11011010", B"00110000",
 B"11011010", B"11011100", B"11010100", B"11010100", B"00111100",
 B"00010100", B"00000111", B"00010101", B"11100100", B"11110000",
 B"00101010", B"00101010", B"00100010", B"00110110", B"11000100",
 B"11100000", B"00100110", B"00100110", B"11100101", B"11110010",
 B"00011010", B"00011011", B"11010111", B"11000101", B"11001101",
 B"00110000", B"11100001", B"11111001", B"11000000", B"00110000",
 B"01000111", B"11100011", B"11010100", B"11010010", B"00100010",
 B"11110111", B"00011010", B"11100100", B"11001001", B"00100101",
 B"11010110", B"11100100", B"00111010", B"11010111", B"00011111",
 B"11100011", B"11101001", B"00010010", B"11010110", B"00001111",
 B"11000100", B"11111010", B"11010100", B"00000110", B"00011111",
 B"11011010", B"11100110", B"00011101", B"11111001", B"11111001",
 B"11010011", B"00101010", B"00100101", B"11101100", B"11011101",
 B"11011000", B"00100000", B"00001110", B"00110111", B"00110000",
 B"11010011", B"11011001", B"00101110", B"11111100", B"00110100",
 B"11001111", B"11010111", B"11010010", B"00011000", B"00111001",
 B"00101011", B"00000100", B"00001110", B"11011011", B"00100111",
 B"11010011", B"00100010", B"11101110", B"11111001", B"00001010",
 B"00001100", B"00010010", B"10111100", B"00010111", B"11101000",
 B"00101010", B"00000010", B"11100101", B"00011011", B"11001101",
 B"00010111", B"11101100", B"11101001", B"00011010", B"11001111",
 B"11100100", B"00110111", B"00100100", B"00011011", B"00100000",
 B"11011000", B"00000100", B"11010011", B"11011110", B"00011101",
 B"01000001", B"00100011", B"00101001", B"11011100", B"11011100",
 B"00011010", B"00100111", B"00001011", B"11011101", B"00100101",
 B"11100011", B"00001010", B"00000001", B"00000110", B"11100100",
 B"00110111", B"11110000", B"00001111", B"11000000", B"11100011",
 B"00000010", B"11010010", B"11100011", B"11101100", B"01000001",
 B"00100000", B"11011100", B"00011010", B"11101001", B"00000001",
 B"11110111", B"00010001", B"11010011", B"11010111", B"11010111",
 B"00100001", B"00111001", B"00100101", B"11010011", B"11100110",
 B"00101001", B"11100010", B"11101111", B"11111110", B"11100011",
 B"00100100", B"00101001", B"10110010", B"00101000", B"00101010",
 B"11001111", B"11110011", B"00101011", B"11000011", B"00100011",
 B"00110010", B"00010110", B"11100001", B"00011101", B"11010010",
 B"00110110", B"11010100", B"11110110", B"00011110", B"00011100",
 B"00100010", B"00101000", B"11100111", B"11011001", B"11101010",
 B"11100010", B"00100100", B"11001000", B"00000110", B"11010110",
 B"11010101", B"00110101", B"00000111", B"11110011", B"00010110",
 B"11001100", B"11011010", B"11100000", B"00100010", B"00011010",
 B"11101111", B"00001110", B"00100100", B"11011010", B"11101011",
 B"11101011", B"11100001", B"11100111", B"00001000", B"11111011",
 B"11100101", B"00101010", B"11101110", B"11011110", B"11001010",
 B"11101001", B"11100000", B"00101001", B"00001100", B"00100011",
 B"11100001", B"00011111", B"11100111", B"00100110", B"11100010",
 B"00110001", B"11010010", B"11001010", B"11100000", B"00010101",
 B"00101110", B"11011100", B"00010110", B"11011100", B"11111100",
 B"00110001", B"11100001", B"00111010", B"00101100", B"11101001",
 B"00011110", B"11111011", B"00111001", B"11011110", B"00000101",
 B"10111111", B"00101100", B"11110111", B"00001110", B"11101010",
 B"00000010", B"00010111", B"11101100", B"00110001", B"00101101",
 B"11100100", B"11001101", B"11101010", B"00000111", B"11010110",
 B"00110100", B"00110000", B"00010010", B"00111010", B"10110100",
 B"11011001", B"11100011", B"00100001", B"00100101", B"11100111",
 B"00111000", B"11101000", B"11011000", B"00001111", B"00101100",
 B"00100111", B"11101000", B"00011110", B"11111000", B"00101001",
 B"11100101", B"00101110", B"00111110", B"00010010", B"11001011",
 B"00001001", B"11100011", B"00110100", B"00100011", B"00011000",
 B"01000001", B"00110110", B"00000011", B"00100110", B"00011001",
 B"00010110", B"00100010", B"00000100", B"00011011", B"11010110",
 B"00100110", B"10111100", B"00001011", B"11011010", B"11001101",
 B"11100010", B"00001110", B"00101101", B"00011001", B"00100001",
 B"10110001", B"11001000", B"11111000", B"11101111", B"00011110",
 B"00011001", B"00100100", B"00000111", B"11010000", B"11010100",
 B"00011000", B"11100001", B"00101011", B"11001010", B"11110011",
 B"11011010", B"00011100", B"00100010", B"11101010", B"00100110",
 B"00100011", B"11100100", B"11100110", B"11000111", B"00000111",
 B"11011011", B"11001011", B"00100110", B"00000011", B"11100011",
 B"11001011", B"11110001", B"11101000", B"11010011", B"11011011",
 B"11110000", B"00111001", B"11101110", B"11101101", B"11010110",
 B"11011010", B"01000000", B"00101101", B"00101110", B"00001101",
 B"01000101", B"00011111", B"00100000", B"00100000", B"00011110",
 B"01000011", B"00010011", B"11001110", B"00101010", B"00110010",
 B"11011000", B"11001010", B"00101111", B"11101000", B"00001000",
 B"00100011", B"11010000", B"11011110", B"11101001", B"11001011",
 B"11100010", B"00001011", B"00110110", B"00001100", B"11001011",
 B"00000000", B"11101110", B"00011101", B"11000100", B"11110011",
 B"00101001", B"00010000", B"11101111", B"11011010", B"11000011",
 B"11011010", B"11110110", B"00011001", B"11011011", B"11011101",
 B"11101000", B"11011001", B"00100100", B"11000010", B"00000010",
 B"11001111", B"11001010", B"11011111", B"11011111", B"00011110",
 B"00011111", B"00011111", B"00000111", B"11010111", B"11110000",
 B"00010100", B"11011001", B"00101000", B"11100111", B"11011000",
 B"00011110", B"00101101", B"00011100", B"00110100", B"11100110",
 B"00010101", B"11100011", B"00000011", B"11010001", B"00011100",
 B"00101011", B"11001110", B"00011001", B"00011100", B"11101010",
 B"11010110", B"00100000", B"00010101", B"00110101", B"11001111",
 B"11100010", B"00001111", B"00101110", B"11101001", B"11001111",
 B"00011011", B"00100011", B"11101011", B"00011000", B"00100111",
 B"11101100", B"11110000", B"00011001", B"00101110", B"00100000",
 B"00011001", B"11011000", B"00101000", B"11011100", B"00101101",
 B"11011111", B"00100001", B"11101010", B"11010100", B"00000001",
 B"11101110", B"11100010", B"11100100", B"11101111", B"11101111",
 B"11110000", B"11110110", B"11100110", B"00010110", B"00011001",
 B"00011110", B"00101111", B"00101110", B"00010101", B"11110011",
 B"00001001", B"00100111", B"11110001", B"11111001", B"00000111",
 B"00011111", B"00101000", B"00110001", B"11010101", B"00000100",
 B"11010100", B"00001000", B"11100000", B"11011111", B"00101110",
 B"00001110", B"00100100", B"11100111", B"00100111", B"11111001",
 B"00011000", B"11100110", B"00101101", B"11011111", B"11001000",
 B"11010101", B"00011001", B"11111011", B"11011010", B"11110011",
 B"00100011", B"11011101", B"00100011", B"11100101", B"11100011",
 B"00101011", B"00101101", B"00100100", B"11110001", B"00100101",
 B"00110110", B"10111110", B"00111010", B"00001001", B"11111001",
 B"11100100", B"00011100", B"00011101", B"11011100", B"11100110",
 B"11111000", B"11011100", B"11011100", B"00100100", B"11001011",
 B"01000011", B"00101011", B"11100010", B"00010100", B"00100011",
 B"11100000", B"11010111", B"11110011", B"11100101", B"00011111",
 B"00100111", B"11101100", B"00100001", B"11100110", B"11010101",
 B"00101111", B"11100110", B"00010011", B"11010001", B"11100111",
 B"00111100", B"00001001", B"10111010", B"00001000", B"00010101",
 B"00111011", B"11110101", B"00100000", B"11111100", B"00110001",
 B"11101110", B"11100000", B"00101011", B"00011010", B"00001111",
 B"00010011", B"11001011", B"11111001", B"00010100", B"00101011",
 B"11100100", B"00110101", B"00110110", B"11100010", B"11111000",
 B"00101111", B"00000111", B"11100101", B"00101000", B"00111000",
 B"00000001", B"00001011", B"11001101", B"11100111", B"00101000",
 B"11010101", B"00010111", B"11101100", B"11100001", B"11100110",
 B"00001100", B"00101011", B"11011011", B"11011000", B"00101010",
 B"00100101", B"00010000", B"00100101", B"11101100", B"11000111",
 B"11010110", B"11001110", B"11110111", B"11101000", B"00011111",
 B"00111010", B"00110000", B"00010100", B"00100010", B"11011001",
 B"00110101", B"00010100", B"11001011", B"00010101", B"00101010",
 B"11001111", B"11010011", B"01001001", B"11011011", B"11101101",
 B"11110010", B"00100110", B"00010001", B"11101101", B"00011101",
 B"00011110", B"00100111", B"00001000", B"00100001", B"00011110",
 B"00000001", B"00100011", B"00010100", B"11011000", B"00011001",
 B"11011100", B"11101011", B"11001101", B"00011000", B"00110100",
 B"00100101", B"11001010", B"11010101", B"11001110", B"11011001",
 B"01000000", B"11010000", B"00101001", B"00011101", B"00001110",
 B"00100001", B"11011111", B"00110110", B"11010000", B"00111000",
 B"11110111", B"00101100", B"11010110", B"11100101", B"00111000",
 B"11011010", B"11110111", B"11011110", B"11011011", B"00001001",
 B"11101011", B"00100010", B"11010100", B"11100000", B"11100111",
 B"00010010", B"00110010", B"00101101", B"11001011", B"11100010",
 B"00100011", B"11110100", B"11011001", B"11010100", B"11011011",
 B"11011001", B"00010110", B"11001111", B"11111101", B"11100010",
 B"00101101", B"00101011", B"11100111", B"11011010", B"11100101",
 B"11010100", B"11111010", B"00001100", B"00100000", B"00001100",
 B"00110100", B"11100111", B"11010001", B"00001110", B"11111100",
 B"00100101", B"11110100", B"11100000", B"00011001", B"00011010",
 B"11110000", B"11110000", B"11100010", B"11111011", B"00100000",
 B"00000111", B"00101010", B"00000110", B"00011111", B"11101000",
 B"00001001", B"11101011", B"11011001", B"00110101", B"01000111",
 B"00101000", B"11101100", B"11010111", B"00011010", B"11100011",
 B"11110011", B"11001100", B"11100100", B"00010110", B"00011011",
 B"11001011", B"11100100", B"00000111", B"00100001", B"11101101",
 B"11000101", B"00010000", B"00110111", B"00011010", B"00001001",
 B"00110000", B"00010011", B"00100101", B"00010010", B"00010001",
 B"00101010", B"00101011", B"11110101", B"00001011", B"11101101",
 B"00010001", B"11001100", B"00011111", B"11101101", B"00100101",
 B"11011111", B"11010111", B"11100001", B"00110100", B"00010111",
 B"11100111", B"00000110", B"01001110", B"11100110", B"11010111",
 B"11011110", B"11101000", B"11011001", B"11000011", B"00011101",
 B"00100011", B"11100100", B"11110010", B"11010111", B"11010110",
 B"11101100", B"11101011", B"00100000", B"00101111", B"11011000",
 B"11111000", B"10101010", B"11100000", B"11100000", B"00011111",
 B"00011101", B"00011011", B"11101001", B"00001111", B"11101110",
 B"00001111", B"11011100", B"00000001", B"11101101", B"00011011",
 B"00010111", B"00010111", B"00001110", B"11101100", B"11101011",
 B"11101001", B"00101110", B"11010010", B"00011110", B"11101001",
 B"11101000", B"00111000", B"00011101", B"01000000", B"11101100",
 B"11011011", B"00111001", B"11010100", B"11001001", B"11100011",
 B"11100011", B"00100010", B"00010011", B"11010100", B"11100111",
 B"00010111", B"00111110", B"11010101", B"11000111", B"11000101",
 B"11011100", B"11100001", B"11000111", B"00101011", B"00010001",
 B"00001110", B"00011100", B"00010011", B"00011011", B"11011001",
 B"00010011", B"00110111", B"11110100", B"11010001", B"00100000",
 B"11001101", B"00011110", B"00100011", B"11001110", B"11101000",
 B"11100110", B"11101101", B"11011011", B"11001111", B"11100110",
 B"11011010", B"00000110", B"00100000", B"11100010", B"00110100",
 B"11011001", B"11001011", B"11101001", B"11010110", B"11011111",
 B"00100010", B"00011000", B"00100111", B"00100101", B"00101100",
 B"00100000", B"00110100", B"00010110", B"00100110", B"00101000",
 B"01000001", B"00001110", B"11100010", B"00001110", B"11100000",
 B"11010100", B"11010110", B"00010100", B"00110111", B"11100001",
 B"00001110", B"11001111", B"11110110", B"00010101", B"11010010",
 B"11011110", B"11010011", B"11100011", B"11100011", B"00101110",
 B"00100101", B"11010101", B"00010000", B"11010000", B"11010101",
 B"10110111", B"11011011", B"11011111", B"00111011", B"11101110",
 B"00101001", B"11100001", B"11001101", B"00110100", B"00001110",
 B"00001110", B"11101100", B"11010110", B"00010100", B"00100010",
 B"11010111", B"11111001", B"00010011", B"00011101", B"11100110",
 B"00010111", B"00101100", B"11101100", B"11111010", B"00010110",
 B"11010110", B"10110011", B"00101101", B"00010001", B"00001110",
 B"00100011", B"11101100", B"11101011", B"11110101", B"11011000",
 B"00011010", B"11011111", B"00110001", B"11011011", B"11010100",
 B"00101000", B"11101011", B"01000011", B"00100110", B"00010011",
 B"11100111", B"00100110", B"11011000", B"00010110", B"00101111",
 B"00001111", B"00101110", B"11100110", B"00101100", B"11110001",
 B"00011111", B"11101001", B"00011011", B"00011001", B"11101111",
 B"11011000", B"00111111", B"00010110", B"11110010", B"11101000",
 B"00100011", B"11100111", B"00100100", B"11001111", B"11100011",
 B"11011000", B"00101000", B"00100010", B"00010001", B"11111100",
 B"11100101", B"00110010", B"11010001", B"11011110", B"11101011",
 B"00001000", B"11100001", B"00011110", B"00010000", B"11001010",
 B"11100001", B"11110011", B"11100100", B"11000111", B"00010101",
 B"11011110", B"11101100", B"11011011", B"11001110", B"00000000",
 B"11011011", B"00010100", B"11011100", B"00101000", B"11101001",
 B"00001111", B"11101110", B"11011000", B"00010001", B"00101001",
 B"00011101", B"00101111", B"11011011", B"00011001", B"00011111",
 B"11011101", B"11100011", B"00100010", B"11011011", B"00100011",
 B"00010011", B"00100110", B"10110110", B"00110001", B"11100000",
 B"00011110", B"00110100", B"11010010", B"00011001", B"00011110",
 B"11101101", B"00000001", B"00110010", B"11100100", B"11011100",
 B"11010101", B"11100100", B"11100101", B"00110110", B"00011000",
 B"00100010", B"00101101", B"00100011", B"00101010", B"11101010",
 B"00101000", B"00010010", B"11101111", B"11010011", B"00001110",
 B"00100000", B"00100001", B"00011100", B"00101001", B"00000101",
 B"01010100", B"00000011", B"00011001", B"00011110", B"00011101",
 B"11100101", B"11100110", B"00111000", B"00011011", B"11101110",
 B"11110011", B"11110110", B"00110010", B"11011000", B"00001111",
 B"11110001", B"11010101", B"00011110", B"00001111", B"11111101",
 B"00101100", B"11010101", B"00100000", B"11011011", B"11010110",
 B"00011010", B"00100111", B"11100001", B"11100010", B"00001110",
 B"11010000", B"00100111", B"11001110", B"11101000", B"00001111",
 B"00010100", B"11001110", B"11001110", B"11110010", B"11010110",
 B"00100110", B"11100110", B"00110110", B"11011010", B"00010110",
 B"11100000", B"11110111", B"11010001", B"00100011", B"00111100",
 B"11010000", B"00100001", B"00100000", B"11100001", B"11101000",
 B"00010110", B"00011001", B"11100101", B"11011010", B"00101100",
 B"11100101", B"01000111", B"00001001", B"11001101", B"00101001",
 B"00100110", B"11010101", B"11101110", B"11110111", B"11011101",
 B"11010101", B"00011101", B"00110001", B"00100101", B"00010101",
 B"11001111", B"11100111", B"11100110", B"00100101", B"00011000",
 B"11111001", B"00011110", B"11100000", B"00001001", B"00000111",
 B"11010111", B"11100011", B"11101010", B"00100011", B"11100000",
 B"00101101", B"00110001", B"11010110", B"11011001", B"11110010",
 B"11101110", B"00100001", B"11010100", B"00100011", B"00100111",
 B"00000110", B"11100101", B"00001100", B"00000010", B"11100010",
 B"11101101", B"00111100", B"00101010", B"00010010", B"11011010",
 B"11001110", B"00011010", B"00111011", B"11010000", B"11011100",
 B"00001110", B"11101011", B"11011110", B"11011000", B"11101010",
 B"00011100", B"11100110", B"11111010", B"11100100", B"10101101",
 B"00110010", B"00110111", B"00010010", B"00101110", B"11100100",
 B"11111110", B"00110100", B"00100111", B"11011100", B"00100111",
 B"00010110", B"11001111", B"11011001", B"00110100", B"00101000",
 B"11111000", B"00101101", B"11010011", B"11001101", B"11000100",
 B"00011111", B"00100101", B"11100011", B"00000100", B"11011011",
 B"00010101", B"11111110", B"11111000", B"00011111", B"00010111",
 B"00100000", B"11000010", B"11011101", B"00010011", B"11010100",
 B"11010011", B"11100101", B"11010011", B"11011010", B"11100010",
 B"11011101", B"11001111", B"00001001", B"00010000", B"00100110",
 B"00011110", B"11010111", B"11110001", B"00100101", B"11011101",
 B"00101011", B"11010101", B"11100111", B"00101010", B"00101011",
 B"11100101", B"00011100", B"11100000", B"11111001", B"11001000",
 B"00100010", B"00010001", B"11110011", B"11011000", B"00110001",
 B"00011110", B"00100111", B"00011110", B"11010111", B"11011101",
 B"11010110", B"00011111", B"11011111", B"11000010", B"11101010",
 B"00011010", B"00001000", B"11000111", B"11010100", B"00011100",
 B"00011011", B"11011000", B"11010011", B"00101011", B"00101100",
 B"11100010", B"11110001", B"00011000", B"11101000", B"11001100",
 B"11011001", B"00100100", B"00111101", B"11100111", B"11100000",
 B"11010110", B"11111010", B"00110101", B"00011001", B"11001000",
 B"00001111", B"11101111", B"00011110", B"11100000", B"00100000",
 B"00100100", B"00000001", B"00010010", B"00100010", B"11010110",
 B"00100010", B"11100011", B"11101100", B"10111100", B"11101001",
 B"00110001", B"11010011", B"11111101", B"00100110", B"00101001",
 B"11101100", B"00111011", B"00010011", B"11001011", B"11100100",
 B"00011111", B"11001110", B"11100010", B"00100011", B"00001111",
 B"00100001", B"00010111", B"11010001", B"11011000", B"11110011",
 B"11100001", B"00011011", B"11101000", B"00011011", B"11100101",
 B"11100100", B"00001110", B"11010100", B"00110001", B"11111010",
 B"00100100", B"11011100", B"00110001", B"11100001", B"00001100",
 B"00100000", B"00110011", B"00011010", B"00101000", B"00001111",
 B"00100101", B"00010101", B"00100001", B"00110001", B"11101011",
 B"11010001", B"00011110", B"11011000", B"11101011", B"11100011",
 B"10111111", B"11011101", B"00001101", B"11101100", B"11110100",
 B"11011010", B"11110100", B"00001110", B"11101100", B"00010110",
 B"00011111", B"11010101", B"11101111", B"00011110", B"00000011",
 B"10110111", B"00000011", B"00100100", B"00011010", B"00101011",
 B"11011011", B"00010101", B"11011100", B"00111001", B"11010110",
 B"11001110", B"11101100", B"11111000", B"11010100", B"00101110",
 B"00001010", B"00100001", B"00110101", B"00011001", B"00100011",
 B"11100010", B"00100100", B"00110011", B"11110011", B"11100101",
 B"00010101", B"11101010", B"11101111", B"00010110", B"11110100",
 B"00111001", B"00001100", B"11101111", B"01000001", B"00100000",
 B"00000110", B"00010100", B"11101011", B"00011110", B"10111110",
 B"00011111", B"11010110", B"00001101", B"11001000", B"00110111",
 B"11001000", B"11100111", B"11011000", B"00110101", B"00011110",
 B"00011101", B"11101110", B"11010011", B"00000011", B"10110001",
 B"00101010", B"11101011", B"00001001", B"11011111", B"00010010",
 B"00010011", B"00100000", B"11001100", B"00010001", B"11100010",
 B"00000101", B"11000000", B"00100100", B"11100011", B"00001101",
 B"10111000", B"11001100", B"00100101", B"00111000", B"00001001",
 B"01010001", B"00010010", B"00000101", B"00101000", B"00110110",
 B"00000111", B"00011111", B"11110011", B"11111011", B"11100000",
 B"00100011", B"01001110", B"11010110", B"00010100", B"11010101",
 B"11011101", B"11010110", B"11110100", B"11010000", B"00100010",
 B"00100010", B"00110001", B"00011110", B"11010110", B"11101010",
 B"11100111", B"11101111", B"00111000", B"00010110", B"00110001",
 B"00010110", B"11000001", B"11010101", B"11011010", B"11100000",
 B"00010000", B"00111010", B"00011010", B"00101111", B"11010010",
 B"00011001", B"11001101", B"11011110", B"11100111", B"00001111",
 B"00001111", B"11100010", B"11001000", B"11011000", B"11100011",
 B"00001010", B"00100111", B"11101100", B"00100010", B"11011100",
 B"11111111", B"00011011", B"11100001", B"11110110", B"11100101",
 B"00011100", B"11111100", B"11110101", B"11010101", B"11101010",
 B"11110110", B"11100111", B"11111101", B"00011100", B"00010000",
 B"00010011", B"00001000", B"00101001", B"00011000", B"11100111",
 B"00010110", B"11100000", B"00011100", B"11100000", B"11100111",
 B"01000010", B"00010111", B"11101100", B"11011111", B"11100101",
 B"11010100", B"11010011", B"00011110", B"00000000", B"00011001",
 B"11110010", B"11110010", B"11010110", B"00101001", B"00100101",
 B"00110101", B"00011011", B"11100111", B"11001100", B"00110101",
 B"00001010", B"11110000", B"10111101", B"00001001", B"00010010",
 B"00011001", B"11011001", B"00110100", B"11011000", B"00001111",
 B"11011100", B"00101110", B"11011110", B"11110001", B"00011110",
 B"11010111", B"11011010", B"11011111", B"11100101", B"11100111",
 B"00100010", B"11110100", B"11110010", B"11011111", B"11111001",
 B"11110010", B"11101011", B"00101101", B"00110010", B"11001011",
 B"00000001", B"00010111", B"11010101", B"11000101", B"00001101",
 B"00011111", B"11011100", B"11011101", B"11001110", B"11100101",
 B"00010111", B"11100010", B"00110000", B"11000100", B"11100011",
 B"11110110", B"11001000", B"00100111", B"00101010", B"00011100",
 B"00011011", B"11011001", B"11001110", B"00100011", B"11011100",
 B"00100010", B"11111111", B"11011101", B"00100011", B"11100110",
 B"11110000", B"11010111", B"00110000", B"00101100", B"11100010",
 B"00100110", B"11001000", B"00010110", B"11011011", B"11010100",
 B"00000110", B"00000011", B"11010101", B"11110010", B"11001100",
 B"11100101", B"00101010", B"11011011", B"00010000", B"11101011",
 B"11100011", B"00101010", B"00101011", B"11011010", B"11001101",
 B"11110000", B"00010100", B"00111111", B"11110000", B"00111011",
 B"11100110", B"11110010", B"11101101", B"00010110", B"00100010",
 B"00001111", B"00101110", B"11100111", B"11101010", B"11010111",
 B"11100001", B"00100100", B"00011000", B"00000101", B"00000011",
 B"11001001", B"11100011", B"11101010", B"11100010", B"11000111",
 B"00101001", B"00100001", B"11110001", B"00010100", B"11111001",
 B"11110111", B"11101101", B"11100101", B"11010001", B"00011111",
 B"00010001", B"00011110", B"00100000", B"00010001", B"00100110",
 B"00110101", B"11010110", B"00000111", B"11011000", B"00101100",
 B"11101110", B"11101011", B"00100110", B"11010100", B"00100000",
 B"11011001", B"11011100", B"00110101", B"01000101", B"00101010",
 B"11100101", B"11111110", B"11010010", B"11100010", B"00010101",
 B"11001000", B"00001110", B"00100111", B"11100011", B"11001000",
 B"11101100", B"10111010", B"00011001", B"11001110", B"00011100",
 B"11011000", B"00101010", B"11011001", B"11100101", B"11101010",
 B"00110101", B"00000011", B"11001001", B"11100011", B"00011101",
 B"00011010", B"00001010", B"11100100", B"00011111", B"11010011",
 B"00011001", B"11101111", B"00100011", B"11000101", B"11011110",
 B"11101010", B"00101011", B"00010100", B"11011111", B"00110010",
 B"00011000", B"00110000", B"00110100", B"00100000", B"00100100",
 B"00111100", B"00001011", B"00011101", B"00001000", B"11110001",
 B"11001010", B"00100111", B"00010001", B"11011001", B"11101110",
 B"00001011", B"11011111", B"00010011", B"00010010", B"11000100",
 B"00001110", B"00111010", B"11010111", B"11001111", B"00101010",
 B"00101110", B"11101010", B"11011100", B"11111100", B"11100010",
 B"11101011", B"00100101", B"11011111", B"11100010", B"00011110",
 B"11100101", B"11011111", B"11010001", B"11101001", B"00101100",
 B"00011010", B"11101101", B"00110101", B"00111011", B"00011010",
 B"11010011", B"00011011", B"11010001", B"00111101", B"00001111",
 B"00100111", B"11001010", B"00100000", B"11011111", B"00101100",
 B"00110001", B"00001100", B"00011110", B"00000011", B"00100101",
 B"11101100", B"00001100", B"11000100", B"11100010", B"11101111",
 B"00101010", B"11001011", B"00100100", B"11001010", B"11001111",
 B"00101010", B"11101010", B"11010110", B"00110111", B"11001100",
 B"00010101", B"11100110", B"11100111", B"00100110", B"11000111",
 B"00100111", B"11011011", B"01001110", B"11100010", B"11101001",
 B"00100010", B"00010111", B"00101111", B"11110000", B"00100110",
 B"11101000", B"00011000", B"11011011", B"00110100", B"11011011",
 B"11100111", B"11100110", B"00100001", B"00100111", B"00110001",
 B"00110010", B"11000011", B"11011011", B"00110010", B"00100110",
 B"00010011", B"00001110", B"00100011", B"00110111", B"11110010",
 B"00011010", B"11100010", B"11001000", B"00110011", B"11011110",
 B"00110000", B"11000011", B"00000010", B"00100001", B"00010100",
 B"00011110", B"11101011", B"00011111", B"00111111", B"10110101",
 B"11110011", B"00011000", B"11110110", B"11010000", B"11111010",
 B"11100010", B"00110101", B"00100110", B"00110010", B"00110111",
 B"11001101", B"00100110", B"00010000", B"11100100", B"11010011",
 B"11101010", B"11000101", B"11001001", B"11001011", B"11111001",
 B"00011010", B"00110010", B"11001001", B"00001101", B"11011000",
 B"00001101", B"00100111", B"11101100", B"00011000", B"01000011",
 B"11110001", B"00110000", B"00010110", B"11101111", B"11010101",
 B"11101001", B"11010110", B"11001001", B"00110011", B"00100001",
 B"00000001", B"00011111", B"00100110", B"11011010", B"11101100",
 B"11010100", B"11011100", B"00100000", B"11110010", B"00011011",
 B"11010101", B"00101010", B"11101100", B"11100101", B"11101000",
 B"00010110", B"00100011", B"11101001", B"00101100", B"11010111",
 B"11011110", B"00010101", B"11000011", B"11010010", B"11001011",
 B"11011011", B"00011100", B"00111011", B"00101100", B"00111001",
 B"00110111", B"00001111", B"00011001", B"00101001", B"00110011",
 B"00111010", B"00001001", B"11111001", B"00101111", B"11001111",
 B"00001010", B"11010111", B"00110011", B"00010000", B"11010000",
 B"00111001", B"00100000", B"11100010", B"11011110", B"00111110",
 B"11011111", B"11110010", B"00010110", B"11100000", B"00010010",
 B"11001011", B"10111010", B"00101001", B"00001100", B"11100010",
 B"11111100", B"11101011", B"11101001", B"11010100", B"11011110",
 B"11101011", B"00011010", B"11001111", B"11111001", B"00001001",
 B"11011011", B"11100100", B"11100111", B"11011111", B"00011010",
 B"11100010", B"00011101", B"11101010", B"11100101", B"11011010",
 B"01000000", B"00011010", B"00000110", B"11101000", B"11001010",
 B"11001111", B"00100000", B"00100000", B"00110101", B"00100010",
 B"00101010", B"00010111", B"11011011", B"11100110", B"00001001",
 B"00110110", B"00000011", B"11101110", B"11011111", B"11011010",
 B"11010010", B"00100101", B"00010101", B"11100000", B"01000000",
 B"11101001", B"00011001", B"11011000", B"00100010", B"11011100",
 B"11010100", B"11100111", B"00101110", B"00010110", B"11101111",
 B"00010101", B"11101111", B"00110010", B"11100001", B"11100101",
 B"00100110", B"00010011", B"11010110", B"00001100", B"00000110",
 B"00100001", B"01000111", B"00110101", B"11100000", B"11100000",
 B"00000011", B"11010010", B"00010110", B"11001101", B"11010111",
 B"11101111", B"00000000", B"00011111", B"11011101", B"11100001",
 B"00111000", B"00011001", B"00101011", B"00101101", B"11100111",
 B"11011111", B"00010011", B"11001101", B"11100010", B"00100010",
 B"11011100", B"11010110", B"11001010", B"11001111", B"00000011",
 B"00011000", B"11101101", B"00001110", B"00011110", B"11101100",
 B"11010100", B"00000011", B"00110010", B"00110110", B"00101001",
 B"11101011", B"00101101", B"11010010", B"00110100", B"11001100",
 B"00000111", B"00101110", B"00110010", B"00011000", B"00101000",
 B"00001101", B"00101010", B"00101000", B"11010100", B"11100101",
 B"01010111", B"11011110", B"00000010", B"11001010", B"11000100",
 B"00001111", B"11101110", B"00101001", B"00101101", B"11100101",
 B"11011010", B"11000111", B"11000101", B"11101101", B"00110100",
 B"00000100", B"00101011", B"11110001", B"00010100", B"11011001",
 B"00100000", B"11101010", B"00101100", B"11011111", B"01000101",
 B"00111101", B"11111100", B"00100011", B"00000110", B"11000000",
 B"11100100", B"11110010", B"11101001", B"00001110", B"00010011",
 B"11010011", B"00011101", B"11001000", B"11000000", B"00101101",
 B"00101011", B"00011011", B"10111010", B"00011011", B"11100101",
 B"00010011", B"00010111", B"11101110", B"11100001", B"00100101",
 B"11100010", B"11100111", B"11101101", B"11001100", B"11001011",
 B"11011101", B"00100101", B"00010010", B"00100010", B"00011010",
 B"11010001", B"11011001", B"11010000", B"00100010", B"00101110",
 B"00010010", B"11011101", B"00110101", B"11011111", B"00001101",
 B"11111001", B"11100100", B"00011000", B"00011011", B"00011110",
 B"00100011", B"11010001", B"11011111", B"00110101", B"11101101",
 B"11100101", B"11100110", B"11100101", B"00110010", B"11101110",
 B"00011011", B"11110011", B"00101101", B"00110000", B"11011001",
 B"11101011", B"11101110", B"11011100", B"11011001", B"11010001",
 B"00010101", B"01000010", B"11101000", B"11000010", B"11010010",
 B"11101101", B"11011011", B"00010110", B"11100010", B"11001001",
 B"00100001", B"11111101", B"00000001", B"11011011", B"11010111",
 B"11100100", B"00010010", B"11100100", B"00001010", B"11101101",
 B"11100110", B"00101011", B"00010110", B"00011001", B"00011111",
 B"00011111", B"11011100", B"00100101", B"11000010", B"00100000",
 B"11100010", B"00001110", B"11100100", B"11001110", B"00010010",
 B"11011111", B"11101110", B"11011000", B"11110101", B"00111011",
 B"00001011", B"00010101", B"11101001", B"00100010", B"11001111",
 B"00101110", B"11100011", B"00100011", B"11001101", B"00110000",
 B"11110010", B"11101000", B"11010001", B"00000110", B"00110011",
 B"11011010", B"00011010", B"00100011", B"00111100", B"10110110",
 B"00100010", B"11100001", B"00000100", B"00001111", B"11001111",
 B"00011001", B"11100111", B"11011011", B"11011100", B"00010101",
 B"00111111", B"00101111", B"11011101", B"00101001", B"11111110",
 B"11011110", B"11101110", B"00110010", B"00101000", B"00001101",
 B"11101010", B"10111101", B"11110100", B"11101101", B"00001111",
 B"11101101", B"00010111", B"00100010", B"00100001", B"00100101",
 B"00101011", B"00101111", B"00110011", B"00001100", B"00010011",
 B"00110001", B"11101101", B"11110100", B"11011100", B"11001101",
 B"00100111", B"11101000", B"00010010", B"11110001", B"11011111",
 B"00111001", B"11001011", B"00010111", B"11011000", B"11100010",
 B"00101000", B"00010110", B"00011100", B"11101011", B"00100100",
 B"00100100", B"11110000", B"11110110", B"00100111", B"00101011",
 B"00010101", B"00101011", B"11100011", B"00110011", B"11100110",
 B"11111010", B"11100001", B"00010011", B"11010001", B"00100111",
 B"00110100", B"11100000", B"00100110", B"00010111", B"11011111",
 B"00100011", B"00010110", B"11000110", B"11010111", B"00100100",
 B"00000111", B"11110011", B"11101011", B"11000110", B"11110000",
 B"11001110", B"00001010", B"00010110", B"11100011", B"01001010",
 B"00000101", B"00100001", B"11101000", B"00010011", B"00100011",
 B"11011000", B"00100000", B"00110010", B"11011100", B"11011100",
 B"11101101", B"11101011", B"00100110", B"00101001", B"11110110",
 B"00001001", B"11000110", B"11101010", B"00100010", B"00110001",
 B"00001100", B"11011100", B"00100101", B"11110011", B"00010001",
 B"00011100", B"11110101", B"11011101", B"00111000", B"11001011",
 B"11110101", B"11001100", B"11101011", B"11011010", B"00101011",
 B"00101110", B"11010111", B"11111001", B"11100000", B"11100111",
 B"11101110", B"11000111", B"11100001", B"00011000", B"11011011",
 B"11111011", B"11001101", B"11000110", B"00000100", B"00101011",
 B"11010111", B"11111100", B"00101111", B"11100101", B"00011010",
 B"00001001", B"11110010", B"00100000", B"11101010", B"11001110",
 B"11010000", B"11100001", B"00100101", B"11100000", B"00101011",
 B"11101111", B"00101001", B"00000000", B"00101010", B"11101001",
 B"01000001", B"11101001", B"00011011", B"11000011", B"00011000",
 B"11011001", B"11010111", B"11000100", B"00011111", B"00010011",
 B"11100010", B"00010000", B"00011010", B"11001101", B"00110000",
 B"00101000", B"11101011", B"11011111", B"00110110", B"00010111",
 B"11101010", B"11111100", B"11100001", B"11010000", B"00010000",
 B"10111001", B"01000110", B"00100011", B"00100101", B"11101001",
 B"00001111", B"00011101", B"11100110", B"11001110", B"00101000",
 B"11101110", B"00101000", B"00101101", B"00010101", B"11100011",
 B"00101001", B"11101010", B"00010011", B"00010000", B"11011110",
 B"11101011", B"00100000", B"11000011", B"11101111", B"11110001",
 B"11010100", B"00101100", B"00101000", B"00010101", B"00101100",
 B"00110101", B"00101001", B"00101100", B"00011001", B"11001011",
 B"00000011", B"00100010", B"00100000", B"11010001", B"00011101",
 B"11111110", B"00110011", B"00000010", B"11100001", B"01001111",
 B"00000101", B"11100000", B"11001011", B"00011010", B"00111101",
 B"11101011", B"11010111", B"00011111", B"11001111", B"00011110",
 B"11011010", B"11000000", B"00110011", B"00111001", B"00001110",
 B"11101111", B"00101100", B"00101111", B"11101010", B"11110011",
 B"00010101", B"11100010", B"11111010", B"00010011", B"00001111",
 B"00110010", B"00001000", B"11100000", B"00000011", B"11011111",
 B"00011101", B"11010110", B"00100111", B"11001101", B"10111000",
 B"00101111", B"00010001", B"00011001", B"00101010", B"00101100",
 B"00111010", B"00011000", B"00010100", B"00010101", B"00100101",
 B"11010001", B"11011100", B"11001101", B"11011111", B"00011011",
 B"00010100", B"11110000", B"00001000", B"11010101", B"00110101",
 B"00111101", B"11011000", B"11111001", B"11001010", B"11011101",
 B"11001000", B"00100011", B"00100010", B"00011010", B"00101000",
 B"00011100", B"00110000", B"00010110", B"00101000", B"11100001",
 B"00010101", B"00010010", B"11011101", B"11101110", B"11110101",
 B"00001011", B"11110101", B"00100101", B"11110100", B"00010101",
 B"11100001", B"11010100", B"11010111", B"00001011", B"00110010",
 B"00010001", B"11101001", B"11011110", B"11000110", B"11011001",
 B"00110000", B"11101110", B"00000110", B"11011110", B"00010011",
 B"00110011", B"00100101", B"11011101", B"00000101", B"11110111",
 B"00001101", B"11100100", B"11111001", B"11101111", B"00011011",
 B"00101001", B"00001111", B"11011001", B"10111011", B"00101000",
 B"00010011", B"11110000", B"00111111", B"00001111", B"11100001",
 B"11001010", B"00100001", B"00001110", B"00010100", B"00010101",
 B"11001001", B"00100111", B"10110111", B"00100000", B"11001111",
 B"00010011", B"00010001", B"11010110", B"00011010", B"00110000",
 B"11010100", B"11011101", B"00001101", B"11000100", B"00101101",
 B"11100010", B"11111011", B"11110000", B"00101010", B"00010010",
 B"10111110", B"11100000", B"00101000", B"00100010", B"00100011",
 B"11110001", B"00000011", B"10111110", B"00001010", B"00010011",
 B"00011101", B"11101000", B"00010001", B"00100111", B"11100001",
 B"00000101", B"00011011", B"00111000", B"00011011", B"00001011",
 B"00011010", B"00100011", B"00010111", B"00011011", B"00101101",
 B"00101000", B"11010100", B"00101101", B"00111000", B"11111001",
 B"00001111", B"00101010", B"11100010", B"00001010", B"00010111",
 B"11010110", B"00011100", B"00100111", B"11111001", B"11101010",
 B"00010011", B"00010111", B"00110101", B"00010010", B"11100010",
 B"00110001", B"11011101", B"00100000", B"11111110", B"00001101",
 B"11011101", B"00101100", B"00101000", B"11011010", B"00011010",
 B"00010111", B"11110001", B"11100100", B"00011011", B"11110101",
 B"11011011", B"11100100", B"00110010", B"00010111", B"11011100",
 B"00100001", B"00010100", B"00101110", B"11101000", B"00110100",
 B"11010100", B"00010010", B"11010100", B"11011000", B"11110111",
 B"00100100", B"00110111", B"00010000", B"00011000", B"11011110",
 B"11100101", B"11100110", B"11000110", B"00101001", B"00010001",
 B"00100100", B"00001110", B"11100011", B"11011001", B"00001000",
 B"11100101", B"11010101", B"00101001", B"11010100", B"11010000",
 B"11011111", B"11001111", B"11010001", B"00100011", B"00000000",
 B"11000110", B"11101011", B"11100011", B"11011011", B"11101000",
 B"00100101", B"11010111", B"00101111", B"00010010", B"11101011",
 B"00100010", B"00110010", B"11010100", B"00101000", B"11101000",
 B"00011000", B"11100110", B"11001010", B"11101000", B"00100010",
 B"00001100", B"11111000", B"11010111", B"11101001", B"00100001",
 B"00000011", B"11111010", B"00101100", B"11001111", B"11011110",
 B"00101011", B"11010010", B"00001000", B"11110100", B"11100000",
 B"00010000", B"00100100", B"00100010", B"00100010", B"00100011",
 B"11011101", B"00100100", B"11010011", B"00100101", B"11011100",
 B"00001101", B"11011010", B"11011000", B"00100100", B"11010111",
 B"11010111", B"11001110", B"11101110", B"00000100", B"11001000",
 B"00001111", B"00000001", B"11110101", B"00011001", B"00110100",
 B"11110011", B"11110010", B"11011010", B"11100001", B"00011010",
 B"00000000", B"11010001", B"00101000", B"11011110", B"00001010",
 B"11100010", B"11100111", B"11110101", B"11101101", B"00011000",
 B"11011111", B"00001011", B"11100100", B"11011110", B"11000101",
 B"11010111", B"00111110", B"01000010", B"00100101", B"00101001",
 B"11101011", B"11011101", B"11101110", B"11111111", B"00011111",
 B"11101011", B"00110000", B"11100010", B"00110011", B"00001001",
 B"00011000", B"11100011", B"00011001", B"11101001", B"00100110",
 B"11011000", B"11100011", B"11011110", B"00001100", B"00101111",
 B"11110011", B"00100010", B"11010011", B"11010011", B"00011010",
 B"11010111", B"00011100", B"11101001", B"11010100", B"10111110",
 B"00011011", B"00110100", B"00100111", B"00010000", B"00101101",
 B"00111000", B"00001011", B"00011100", B"00100101", B"00111000",
 B"11100001", B"11010001", B"00100100", B"00100100", B"00001101",
 B"00111011", B"11111001", B"11100010", B"00011110", B"00100111",
 B"11011010", B"11101001", B"00011011", B"00101000", B"11101001",
 B"11110001", B"11110001", B"00000110", B"00000110", B"11001101",
 B"11001111", B"11101111", B"11101110", B"11100000", B"00100111",
 B"11001110", B"00011001", B"11101100", B"11011101", B"11110001",
 B"00101001", B"00011001", B"00001110", B"11110000", B"00110011",
 B"11011110", B"11011000", B"11101000", B"00000000", B"00110001",
 B"11101010", B"11011000", B"00100001", B"00100001", B"00101101",
 B"00110111", B"11110110", B"11001011", B"00110000", B"00101011",
 B"00011011", B"01000100", B"00101010", B"00011101", B"00100011",
 B"00010110", B"01001101", B"11000111", B"00011000", B"00101110",
 B"11010101", B"00001011", B"00010000", B"11101000", B"11101000",
 B"00011001", B"11100110", B"11100110", B"11010011", B"00101101",
 B"00100010", B"11100000", B"11011111", B"00001111", B"11101000",
 B"11100111", B"11101111", B"00011101", B"00011010", B"11111100",
 B"00111110", B"01000010", B"00000010", B"11010011", B"00100100",
 B"11011001", B"00011001", B"11100011", B"11011011", B"00101000",
 B"11111000", B"11011101", B"11011111", B"00100000", B"00110000",
 B"11011101", B"11100010", B"00100010", B"00110000", B"11101010",
 B"11100111", B"11100110", B"11100000", B"11100001", B"11000010",
 B"11100000", B"11001001", B"11001000", B"00011110", B"00100110",
 B"00110010", B"00011000", B"00100011", B"11100000", B"00000100",
 B"00011101", B"11110100", B"00100110", B"00011111", B"11101101",
 B"11101100", B"00011101", B"00011000", B"11100101", B"11111001",
 B"11100000", B"11011101", B"11101001", B"00011011", B"00011010",
 B"00001110", B"11100011", B"00001011", B"00100010", B"11100010",
 B"11100000", B"00111010", B"00001000", B"00101110", B"00010000",
 B"00100100", B"00011111", B"00001101", B"00011111", B"11001100",
 B"00011110", B"11100000", B"00011111", B"11011011", B"00000111",
 B"00010000", B"00100000", B"11101000", B"00101011", B"00101101",
 B"00010110", B"11001101", B"00101000", B"11011110", B"00011100",
 B"00011000", B"11010110", B"10111011", B"00101110", B"11110010",
 B"11011100", B"11011100", B"11011110", B"11001100", B"00011100",
 B"01000111", B"00110010", B"11011110", B"00101000", B"11101111",
 B"00011000", B"00110011", B"00100100", B"00000001", B"00101011",
 B"00110111", B"00100001", B"00010011", B"00101001", B"11011001",
 B"11110011", B"00010000", B"11010000", B"00100101", B"11010101",
 B"11011111", B"00100100", B"00100100", B"11100101", B"00011111",
 B"00100110", B"11100100", B"00100101", B"00000111", B"11011001",
 B"11101110", B"11100000", B"00110010", B"00110110", B"00101001",
 B"00011010", B"11110001", B"11001010", B"11100010", B"11011001",
 B"11101110", B"00010110", B"00110011", B"11010011", B"00011101",
 B"11111110", B"00011111", B"00101000", B"00011000", B"11000111",
 B"00001001", B"11110000", B"00011010", B"11101101", B"00101100",
 B"11110000", B"11101101", B"11010011", B"11100111", B"00101001",
 B"11011101", B"11111011", B"00010100", B"00100101", B"00010101",
 B"11100100", B"00100001", B"11000011", B"00111001", B"11010010",
 B"00100010", B"11000000", B"00100010", B"11101001", B"11100100",
 B"11101000", B"00010011", B"00010011", B"00100000", B"00010111",
 B"00100011", B"11001011", B"00101000", B"11110000", B"00100010",
 B"11011000", B"00010110", B"11110000", B"00101000", B"11101101",
 B"11110010", B"11100000", B"00010011", B"11111011", B"11011100",
 B"00110111", B"00110101", B"00100000", B"11101010", B"00011100",
 B"11111101", B"00100001", B"11001101", B"11111111", B"11001111",
 B"11010111", B"00101001", B"00011001", B"00100111", B"00101000",
 B"11100101", B"00011101", B"00110111", B"00100000", B"11100111",
 B"00100101", B"11001110", B"01001000", B"00010010", B"11101010",
 B"11110001", B"11101111", B"11011101", B"00100000", B"11100000",
 B"00100100", B"11110110", B"11100001", B"00011011", B"00100001",
 B"00011011", B"00010001", B"11010001", B"11011110", B"00001001",
 B"11010101", B"11011011", B"11001110", B"11011100", B"00100000",
 B"11110000", B"00011110", B"11010101", B"00101010", B"11011100",
 B"00011100", B"11101010", B"11001111", B"00100101", B"00000100",
 B"00011101", B"00011101", B"11111010", B"11101100", B"00110101",
 B"00001101", B"11010101", B"11100011", B"11111110", B"00001101",
 B"11011100", B"00100000", B"00001000", B"11011011", B"11100011",
 B"00110000", B"00001000", B"11110110", B"00101001", B"11110110",
 B"00100000", B"11011111", B"11100001", B"00011100", B"00111110",
 B"00010101", B"11110111", B"11011111", B"00010010", B"00011111",
 B"11111001", B"11110001", B"11111000", B"00100101", B"11100100",
 B"11010101", B"11011000", B"00110110", B"00101000", B"11001010",
 B"00100001", B"11100001", B"00001101", B"00110011", B"11100100",
 B"00101001", B"01000111", B"11010111", B"11100010", B"11010101",
 B"11111000", B"11101001", B"00100010", B"00101000", B"00110101",
 B"00100110", B"00010000", B"11101011", B"00110101", B"10110110",
 B"00011000", B"11000000", B"11001100", B"00111011", B"11010001",
 B"11110101", B"00001101", B"00001001", B"00011010", B"00011000",
 B"11100001", B"11100011", B"11011111", B"00111100", B"00010110",
 B"00101000", B"11111110", B"00101011", B"11011100", B"00100111",
 B"00100010", B"11010110", B"11111111", B"00100111", B"11011011",
 B"00100100", B"00010011", B"11101001", B"11100100", B"00111000",
 B"00101011", B"11111001", B"11010100", B"11100101", B"11011111",
 B"11010001", B"00011110", B"00001101", B"11110101", B"11100111",
 B"00011100", B"00011000", B"11011000", B"11100000", B"11010101",
 B"11011010", B"11010001", B"00011010", B"00011010", B"11100110",
 B"00010111", B"11110010", B"00100010", B"10111100", B"00100011",
 B"11011111", B"11011000", B"11011011", B"00001100", B"00011011",
 B"00011101", B"11100111", B"00001001", B"11001100", B"11100010",
 B"11111101", B"00111110", B"00001100", B"11000010", B"10111001",
 B"00100001", B"00011100", B"00110101", B"00011001", B"11011010",
 B"00000011", B"11011011", B"11000101", B"11011111", B"11100011",
 B"00101011", B"00110011", B"00101110", B"00111111", B"11111000",
 B"11011111", B"00011110", B"00011101", B"00011100", B"00100101",
 B"11000101", B"11101110", B"11100000", B"11101101", B"00011101",
 B"00100000", B"00011010", B"00100000", B"11101001", B"11001110",
 B"00100010", B"00010011", B"00010111", B"11001111", B"00011100",
 B"11011101", B"11111001", B"11010010", B"11110000", B"11101000",
 B"11101011", B"00011110", B"00001101", B"11101101", B"00110110",
 B"11101100", B"11101001", B"00101001", B"00001110", B"00000111",
 B"11011000", B"00011101", B"11100111", B"00100010", B"00001100",
 B"11010010", B"00001100", B"11110100", B"11100010", B"11100110",
 B"00100101", B"00101011", B"11101110", B"11011101", B"11110001",
 B"11001011", B"00100010", B"00001111", B"00111001", B"00010101",
 B"00110011", B"11110101", B"00100001", B"11100111", B"11100001",
 B"11011010", B"00011000", B"00010110", B"11010111", B"00100010",
 B"11011011", B"11001101", B"11001011", B"00010110", B"00110000",
 B"11000100", B"11100100", B"11010001", B"00011100", B"11011110",
 B"00100101", B"11101000", B"11000010", B"00011000", B"11011111",
 B"00100010", B"00001100", B"11100011", B"11010100", B"11100000",
 B"11100011", B"11101100", B"11011011", B"00011101", B"11011111",
 B"10110111", B"11011011", B"00100000", B"00100000", B"11101000",
 B"11100101", B"11100111", B"11010100", B"11101010", B"00010000",
 B"00101101", B"01000011", B"00011111", B"00010111", B"00100011",
 B"00011011", B"11100101", B"00101010", B"11001110", B"00010100",
 B"11110011", B"00001111", B"10111100", B"00110000", B"11010111",
 B"11011110", B"11101011", B"00110000", B"00010111", B"00010100",
 B"00111011", B"00010101", B"11010001", B"00100100", B"11111100",
 B"00100101", B"11000100", B"11110100", B"00000011", B"00010110",
 B"00100100", B"11010011", B"00000101", B"11100110", B"00010110",
 B"11100001", B"11111001", B"00110100", B"00100111", B"00010011",
 B"00110111", B"11011101", B"11101111", B"00110110", B"11001010",
 B"11101100", B"00111101", B"11001110", B"11110011", B"11101010",
 B"11010001", B"11011100", B"00100110", B"11011100", B"00111111",
 B"11100100", B"11100100", B"00111000", B"00100101", B"11001110",
 B"00100011", B"00010010", B"00011100", B"11001110", B"00100010",
 B"00000110", B"00010110", B"00000010", B"00100011", B"11011001",
 B"11110110", B"00010110", B"00110100", B"11011001", B"11100001",
 B"11010001", B"11110000", B"11011000", B"11100101", B"00100110",
 B"00001010", B"00100110", B"00101100", B"00101111", B"00011011",
 B"11001010", B"11100011", B"00101100", B"00010010", B"11100100",
 B"11100011", B"11110001", B"11010111", B"00011001", B"00101110",
 B"00010100", B"00101001", B"11011011", B"11000111", B"11100000",
 B"11011011", B"00011010", B"11011010", B"00010010", B"11010110",
 B"11011001", B"00101000", B"11101000", B"11010111", B"00101110",
 B"11100111", B"00111001", B"11101001", B"11010111", B"00011010",
 B"10111101", B"00011100", B"11000111", B"11100000", B"11100010",
 B"00100011", B"00110010", B"11110000", B"11111000", B"00100011",
 B"00010001", B"00100000", B"00010100", B"00000100", B"00100011",
 B"00101001", B"00111001", B"00110000", B"11101011", B"11100110",
 B"00101110", B"00101110", B"11111100", B"11011101", B"11011100",
 B"00011101", B"00100101", B"00011101", B"11011101", B"00011110",
 B"11100011", B"00111001", B"00011110", B"00100001", B"00010000",
 B"11111010", B"00100001", B"11100001", B"00010010", B"11101011",
 B"00000101", B"00100111", B"11010100", B"11101101", B"00101111",
 B"00101011", B"11010011", B"11110000", B"11100111", B"00100100",
 B"11010110", B"00100111", B"11101010", B"11100111", B"00010100",
 B"00100010", B"11001111", B"00110010", B"00110110", B"00110100",
 B"11100001", B"00111000", B"11110011", B"11111100", B"01010000",
 B"00100111", B"00011010", B"00010101", B"00010011", B"00100100",
 B"00001110", B"00110100", B"00101111", B"00100101", B"00000111",
 B"00110001", B"00101000", B"00010101", B"00100101", B"00011101",
 B"00010010", B"11001011", B"11100010", B"11011000", B"11011011",
 B"00000100", B"11101001", B"00010110", B"11100001", B"11101000",
 B"00000110", B"11100001", B"00010111", B"11100000", B"11100101",
 B"00110100", B"11001001", B"11011010", B"00100111", B"00100111",
 B"00111001", B"00111000", B"11011010", B"11000001", B"10111111",
 B"11011001", B"11100001", B"00010101", B"00101000", B"11100011",
 B"00010011", B"11101111", B"11101101", B"11011010", B"11101000",
 B"11101001", B"00011111", B"00100111", B"00011110", B"00110100",
 B"00010000", B"00100010", B"11100001", B"00101101", B"00101011",
 B"11011001", B"11100110", B"00111010", B"00111000", B"11001100",
 B"11111001", B"00001001", B"11001001", B"00001101", B"00101000",
 B"11101111", B"11010000", B"11100111", B"00101010", B"11010100",
 B"00101110", B"11011010", B"11001010", B"00100110", B"11011111",
 B"00111000", B"00001111", B"00011110", B"11100100", B"00010001",
 B"11100011", B"00010011", B"11110101", B"00001010", B"11010111",
 B"00010110", B"11100101", B"11011010", B"00010011", B"00100011",
 B"11011000", B"00001110", B"11110101", B"11011111", B"11110001",
 B"00110001", B"00110111", B"11011100", B"11101011", B"00101011",
 B"00110100", B"11100010", B"11100011", B"11100110", B"11101111",
 B"11010011", B"00101100", B"00100000", B"11101001", B"00011001",
 B"01000000", B"11010110", B"11100001", B"00011100", B"11001110",
 B"11011100", B"11011111", B"11011011", B"00100110", B"00011110",
 B"00100111", B"00010100", B"11101111", B"00011010", B"11011010",
 B"11101100", B"11101001", B"00101111", B"00100111", B"11110010",
 B"00011101", B"11100111", B"11011011", B"11011111", B"11101000",
 B"00101001", B"11000000", B"00001001", B"11110100", B"00110111",
 B"11010110", B"00011000", B"11011110", B"11100101", B"00011010",
 B"00111111", B"11100001", B"00011011", B"00100000", B"11101001",
 B"11011111", B"11000010", B"11100000", B"11001010", B"11011011",
 B"11101100", B"11101000", B"00101001", B"00011110", B"11010111",
 B"00010001", B"11001111", B"11100100", B"11010110", B"11100111",
 B"00101000", B"00110010", B"11011001", B"00011111", B"11101101",
 B"00100011", B"11001101", B"11011110", B"00001001", B"11011011",
 B"11001110", B"11001111", B"10111001", B"11110010", B"11010111",
 B"00101000", B"11011011", B"00011001", B"11101010", B"11100100",
 B"00010111", B"11110000", B"00011010", B"00010011", B"11001001",
 B"11110010", B"11110100", B"11100011", B"11010111", B"00101011",
 B"11011000", B"00100001", B"11100101", B"11001001", B"11011111",
 B"00110111", B"00101001", B"00010000", B"11010111", B"00010011",
 B"11011000", B"11010010", B"11110010", B"00100111", B"00101100",
 B"11101101", B"11100010", B"00010110", B"11101010", B"00100110",
 B"11011101", B"11010010", B"00101000", B"00000011", B"00010100",
 B"00011011", B"11101111", B"11110110", B"11010101", B"11010100",
 B"11100001", B"00111001", B"11100110", B"00011011", B"11100111",
 B"11101111", B"11110001", B"00010011", B"00001110", B"00011101",
 B"00001011", B"11110100", B"11010000", B"00101000", B"00101110",
 B"11011000", B"11101111", B"11110100", B"00001110", B"00010000",
 B"11010111", B"11100101", B"00100101", B"11101010", B"11101001",
 B"00100100", B"11101101", B"00110000", B"11110011", B"11100000",
 B"11100111", B"00100110", B"00010000", B"00010001", B"11000001",
 B"11001010", B"00010001", B"11101101", B"11101000", B"11110010",
 B"11100111", B"11101110", B"11010110", B"11010001", B"11101100",
 B"00011100", B"00011111", B"00011110", B"00010001", B"11101100",
 B"11011110", B"00100101", B"11110111", B"00100010", B"11101010",
 B"11010000", B"00110100", B"00010001", B"11111001", B"00001110",
 B"00000100", B"11100000", B"00000110", B"00011011", B"11010111",
 B"11110111", B"11011110", B"11011010", B"10111110", B"00000100",
 B"00110001", B"00101101", B"01001100", B"11101110", B"00100100",
 B"11101100", B"11100111", B"11010010", B"00011110", B"00100001",
 B"11110000", B"11100000", B"00110000", B"00100010", B"11010110",
 B"11010010", B"11101110", B"11110101", B"11010001", B"11110101",
 B"00101100", B"00101011", B"10110000", B"11101010", B"00000001",
 B"11100011", B"11101010", B"00010111", B"11010110", B"00001000",
 B"11110100", B"11001110", B"00101011", B"11100010", B"00000011",
 B"11011001", B"00101001", B"00000011", B"00100000", B"11001101",
 B"10111110", B"00100101", B"00111011", B"00011111", B"11110000",
 B"00101110", B"11100001", B"11100111", B"11011111", B"00100101",
 B"00100110", B"00011101", B"00101101", B"11000001", B"00001110",
 B"00100101", B"11101001", B"11110011", B"00011010", B"11010101",
 B"00001010", B"00000101", B"00100011", B"11101101", B"00011101",
 B"11011111", B"11111100", B"11010011", B"00100011", B"11010101",
 B"11001111", B"11100010", B"00100111", B"00100001", B"11101011",
 B"00100101", B"11100110", B"00011101", B"00010001", B"11010011",
 B"00110000", B"00000100", B"11100001", B"00100000", B"11000010",
 B"11011111", B"11100111", B"11011011", B"00110111", B"11010111",
 B"00000100", B"00010101", B"00101010", B"11110101", B"11101000",
 B"00000000", B"00101100", B"11011011", B"11010000", B"11101000",
 B"11011101", B"00000110", B"11001110", B"00110000", B"11011001",
 B"11010110", B"00000100", B"11010001", B"00000011", B"11010100",
 B"11111111", B"00100110", B"00000111", B"00101101", B"11111011",
 B"00100111", B"00011101", B"00010101", B"11011101", B"00000111",
 B"11010111", B"00100110", B"11101001", B"00001111", B"11000001",
 B"00010000", B"11100010", B"11100101", B"10110110", B"00101110",
 B"00100010", B"00001111", B"00011100", B"11010111", B"11010011",
 B"00111011", B"00100011", B"11000000", B"11101100", B"11100110",
 B"11110100", B"00100111", B"00011100", B"11011000", B"00010001",
 B"11101110", B"00010010", B"11101111", B"11010111", B"00011010",
 B"11110000", B"00010101", B"11101100", B"11010001", B"00011101",
 B"00001111", B"00100010", B"00110011", B"11100110", B"00010010",
 B"11100010", B"00101100", B"11010101", B"00100100", B"00100110",
 B"00001001", B"00101000", B"00100000", B"00011110", B"00100001",
 B"00101101", B"00110110", B"11010000", B"11100000", B"11010010",
 B"11100011", B"00100100", B"11011010", B"00100101", B"11100010",
 B"00001101", B"11101110", B"00000110", B"11100100", B"11100100",
 B"01000000", B"00000101", B"11100001", B"00101001", B"00011110",
 B"00011001", B"11010100", B"00100110", B"11100001", B"00001111",
 B"00010111", B"00100111", B"11001101", B"00100011", B"01001101",
 B"11101010", B"11100010", B"00011010", B"00011101", B"00101000",
 B"00100101", B"00010011", B"00101001", B"00111001", B"00101010",
 B"00000010", B"00101101", B"00001001", B"11010000", B"11000100",
 B"00100110", B"00101010", B"11010010", B"11110110", B"00001010",
 B"11100101", B"00011000", B"00010111", B"11101001", B"00101100",
 B"00010111", B"11001111", B"00001011", B"11100100", B"00110000",
 B"00011111", B"11011010", B"00101001", B"00100001", B"11100001",
 B"00111010", B"00100111", B"00110101", B"00100011", B"11111110",
 B"00101101", B"00010111", B"00011110", B"00110011", B"11001000",
 B"11101001", B"11001110", B"11100000", B"00110001", B"11011111",
 B"00100101", B"11101101", B"00010111", B"00001101", B"00101011",
 B"11101001", B"00001111", B"11110010", B"00001101", B"00011100",
 B"11011111", B"00011011", B"11100100", B"11010001", B"11011100",
 B"00010111", B"00010011", B"11001110", B"00110001", B"00011101",
 B"11011111", B"11100011", B"11100111", B"11010111", B"11101011",
 B"11110010", B"11101100", B"11010111", B"11101001", B"00110110",
 B"00010000", B"00001110", B"00011110", B"11001111", B"11100011",
 B"11110101", B"00101100", B"00100001", B"11100100", B"00010001",
 B"11010000", B"00010001", B"00000111", B"11100000", B"00110100",
 B"00001001", B"11010111", B"11010011", B"00110101", B"00011111",
 B"00010100", B"11011100", B"00011010", B"00011100", B"11000010",
 B"11101110", B"01001001", B"00110000", B"00001011", B"00011000",
 B"00011001", B"00011111", B"00111101", B"00010001", B"00011100",
 B"11000100", B"11101000", B"00110011", B"00101001", B"00100001",
 B"00100111", B"11010001", B"11100000", B"00100010", B"00101111",
 B"11001101", B"00010110", B"00101011", B"11100011", B"11001000",
 B"00000001", B"00101011", B"11000101", B"11001000", B"11010001",
 B"11011111", B"00100101", B"11100010", B"00101100", B"00111111",
 B"01000000", B"00100001", B"00101001", B"01000111", B"00010100",
 B"00000100", B"00010101", B"11011110", B"00000000", B"11101011",
 B"11101000", B"11101010", B"00010000", B"00011111", B"11010010",
 B"11100101", B"11011010", B"11010001", B"00101110", B"00011101",
 B"11101101", B"00011111", B"11101001", B"11010111", B"11010000",
 B"00100110", B"11110100", B"00100101", B"00000111", B"11101101",
 B"00110001", B"11101001", B"11011011", B"11001001", B"00001100",
 B"00000101", B"11001010", B"00100111", B"11010111", B"00100111",
 B"00011000", B"00101110", B"00011110", B"00101100", B"00011010",
 B"00010110", B"00101110", B"00110100", B"00010000", B"11110110",
 B"00101111", B"00100001", B"11101101", B"11010001", B"00011100",
 B"11000110", B"00011011", B"00011110", B"11010010", B"11111010",
 B"00000101", B"11001010", B"11011010", B"00101000", B"00011011",
 B"11100101", B"11100001", B"11111101", B"00100111", B"11100000",
 B"11100100", B"11110110", B"11101101", B"11010111", B"11011110",
 B"00011100", B"00111101", B"00011000", B"00010111", B"11101011",
 B"11101111", B"00001110", B"00010111", B"00100100", B"00100001",
 B"11101001", B"11011101", B"00100100", B"00111001", B"00011111",
 B"00101111", B"00000010", B"00100001", B"00011110", B"00110000",
 B"00100100", B"11100100", B"00000100", B"11011000", B"11000111",
 B"11100011", B"00101100", B"11111001", B"11101000", B"11011111",
 B"00111010", B"11001111", B"00000011", B"11100100", B"11000110",
 B"01000010", B"11111010", B"00110111", B"00011101", B"11010101",
 B"00010011", B"11000111", B"00011011", B"11101110", B"11100011",
 B"11001010", B"11111000", B"00011100", B"00100111", B"11100000",
 B"00011001", B"11001110", B"00110101", B"00110011", B"00100000",
 B"11101110", B"00100001", B"11011111", B"00100011", B"11010110",
 B"11010101", B"11100000", B"00010010", B"11101001", B"00101100",
 B"11110111", B"11101000", B"00001001", B"00001101", B"00011100",
 B"00100100", B"00000101", B"00110010", B"00000111", B"00001010",
 B"00011100", B"00011101", B"00101001", B"11011010", B"00011100",
 B"00001100", B"11010010", B"11100000", B"00000001", B"00101011",
 B"11010010", B"11010100", B"00011010", B"11011000", B"11100000",
 B"11100101", B"11010001", B"00000100", B"00010011", B"00000011",
 B"00001100", B"00000111", B"00100001", B"11111110", B"00011011",
 B"00101000", B"00100011", B"11010100", B"00010011", B"00000000",
 B"11101000", B"11010110", B"00101101", B"00011100", B"00001111",
 B"11010001", B"11011011", B"00011001", B"11111110", B"11101000",
 B"11101110", B"00011001", B"11110010", B"00111000", B"00011101",
 B"11110110", B"00011101", B"00100110", B"11010111", B"11111001",
 B"00011110", B"00110000", B"00011000", B"11101100", B"00110000",
 B"11011010", B"00100100", B"11010100", B"00100101", B"11100000",
 B"11100011", B"11101000", B"11111100", B"00011100", B"11001010",
 B"00011001", B"00011001", B"00011011", B"11101000", B"00110010",
 B"11101011", B"00101110", B"11010101", B"11101011", B"11001110",
 B"00010011", B"11110011", B"00100100", B"11001001", B"11100111",
 B"00100101", B"10111101", B"11001101", B"11010100", B"00111010",
 B"00100101", B"11101000", B"00011010", B"11101000", B"11101101",
 B"01000100", B"00101000", B"00101100", B"11010111", B"00011101",
 B"11000001", B"00101111", B"00011100", B"00101001", B"00101001",
 B"11010001", B"00111010", B"11010110", B"00001011", B"11001101",
 B"00011110", B"00110000", B"11110110", B"11101000", B"00011101",
 B"00001011", B"11101101", B"11101111", B"01000111", B"11110000",
 B"00100110", B"00011011", B"11100010", B"00011110", B"00100000",
 B"11100100", B"11010100", B"00011010", B"00111110", B"11110110",
 B"11001100", B"11101010", B"11011001", B"11011011", B"00011101",
 B"11101001", B"00011000", B"11100100", B"11011011", B"11010110",
 B"00100100", B"00100000", B"11011111", B"00101010", B"00011000",
 B"11100011", B"11100011", B"11011100", B"11000100", B"11101000",
 B"00011001", B"00010001", B"11110000", B"00001010", B"00101000",
 B"11110001", B"11010111", B"00010101", B"11110010", B"00011110",
 B"11011010", B"00011000", B"11101010", B"11100010", B"00010000",
 B"00111000", B"00100101", B"01000000", B"00000110", B"11011010",
 B"00110001", B"11011001", B"00101001", B"11011101", B"00010101",
 B"00100010", B"00101111", B"00100000", B"00100110", B"00110111",
 B"00100101", B"00001111", B"11010111", B"00011110", B"11010010",
 B"00011011", B"00000010", B"11110110", B"00101001", B"00100011",
 B"11100111", B"11011001", B"00000011", B"00110100", B"01000000",
 B"11100111", B"00110101", B"11100010", B"00110001", B"11011000",
 B"11101111", B"11110110", B"11101000", B"00100000", B"11111111",
 B"00011110", B"11110101", B"11011011", B"00010010", B"11100000",
 B"00110000", B"11100010", B"11011101", B"00011011", B"11110100",
 B"11110010", B"11100000", B"11011110", B"00000100", B"00011111",
 B"00011001", B"00011000", B"11110010", B"11010010", B"11100001",
 B"11000101", B"00010000", B"11111011", B"00001000", B"01001011",
 B"00110000", B"11011111", B"00100001", B"00101011", B"11110101",
 B"00101001", B"00100100", B"11111000", B"00001001", B"11110101",
 B"11111001", B"11001101", B"00110001", B"00100101", B"00010101",
 B"00101011", B"11010111", B"11011111", B"00110111", B"11010011",
 B"00010011", B"11100010", B"11101001", B"00100001", B"11100111",
 B"11111110", B"11110100", B"00011110", B"00101100", B"11010110",
 B"00101010", B"11100010", B"00001110", B"11010010", B"00001100",
 B"11010101", B"11011100", B"11011101", B"00010010", B"00100011",
 B"00100100", B"11100111", B"11001001", B"11011011", B"11100110",
 B"00011101", B"11100110", B"00011000", B"00100011", B"00011110",
 B"11010101", B"11100001", B"00010100", B"00010101", B"11111110",
 B"11110000", B"11011011", B"11010101", B"00100111", B"11000010",
 B"00011000", B"11100100", B"11011111", B"00101010", B"11011100",
 B"11111000", B"00100101", B"00101011", B"00100010", B"00111100",
 B"11010110", B"00000101", B"11001100", B"00011010", B"11100110",
 B"11011100", B"11101101", B"00001101", B"00010110", B"11101110",
 B"11011110", B"11010100", B"10111100", B"00100110", B"00110100",
 B"10111110", B"00101000", B"11111001", B"11100010", B"11111001",
 B"11111010", B"00001100", B"00110001", B"11100000", B"00011000",
 B"11100111", B"00101100", B"00011100", B"00011111", B"11011101",
 B"00011110", B"11000000", B"00101101", B"11001001", B"00011111",
 B"11010101", B"00111101", B"11011010", B"11011011", B"11011101",
 B"00100010", B"11110111", B"11011100", B"11010000", B"11001010",
 B"00011010", B"00111110", B"11010000", B"00101010", B"11100101",
 B"11010001", B"00011011", B"00101111", B"00101111", B"11101100",
 B"00011000", B"11100000", B"00010100", B"00011000", B"11011100",
 B"11001111", B"11011110", B"11010011", B"00010111", B"11100000",
 B"00110010", B"00011011", B"00010011", B"11010001", B"00011110",
 B"00011011", B"11110000", B"11000101", B"00101001", B"00111000",
 B"11101101", B"11010101", B"00101101", B"11011100", B"11001001",
 B"11101011", B"11011100", B"00001101", B"11101111", B"10110111",
 B"00000101", B"11110000", B"00101100", B"11001110", B"00010110",
 B"11101111", B"00011111", B"11100010", B"11011100", B"11100110",
 B"00010010", B"00101101", B"11011110", B"00010010", B"11010010",
 B"00001100", B"00101001", B"11011101", B"00101001", B"00011110",
 B"11110101", B"11011011", B"11100101", B"11111111", B"00011100",
 B"00101000", B"11001111", B"00101011", B"11110110", B"00010010",
 B"00010111", B"11011110", B"00001100", B"00011001", B"11100001",
 B"11010111", B"00000111", B"00011110", B"00101100", B"00001111",
 B"11001010", B"00011100", B"11100001", B"00101001", B"11011100",
 B"11010110", B"11100100", B"11101110", B"00100000", B"00000101",
 B"11001101", B"00101101", B"11011110", B"00011100", B"11100000",
 B"11001011", B"00011111", B"11011001", B"11010101", B"11111111",
 B"11111100", B"11100111", B"00101100", B"11001110", B"00010100",
 B"11010100", B"11010000", B"00101011", B"00100011", B"00101001",
 B"11101000", B"00111010", B"00000010", B"11011100", B"11110111",
 B"00010000", B"00101001", B"11101010", B"00001010", B"00001100",
 B"00101110", B"11100111", B"00010101", B"11101000", B"00010000",
 B"00100110", B"11100111", B"11100010", B"00101011", B"00000011",
 B"11011010", B"11101010", B"11111001", B"11101101", B"00010010",
 B"11011001", B"00101011", B"11010010", B"11110011", B"00001011",
 B"00101110", B"00101100", B"11100110", B"00100001", B"11110011",
 B"11110010", B"11110000", B"00011010", B"00101011", B"11010000",
 B"11100011", B"00100100", B"00010111", B"00011001", B"00110100",
 B"11100001", B"11010111", B"00001101", B"01000110", B"00011000",
 B"11101011", B"00011001", B"11010111", B"00010100", B"11110100",
 B"11010110", B"00001011", B"00110010", B"11011101", B"11010100",
 B"11011001", B"11001010", B"11101000", B"11100011", B"11001100",
 B"00000001", B"00001100", B"00010010", B"11101100", B"00000000",
 B"11110010", B"11010011", B"00110101", B"00011101", B"00001010",
 B"11001101", B"00010110", B"11101111", B"00111010", B"11110101",
 B"00100101", B"00001011", B"00110001", B"11110001", B"00111010",
 B"11101111", B"00101010", B"11010000", B"11101001", B"11001111",
 B"00110101", B"00011010", B"11110110", B"00110000", B"11000111",
 B"00110001", B"11000010", B"01000001", B"11011101", B"11100100",
 B"11110101", B"00001001", B"00100110", B"00101111", B"11110110",
 B"00101010", B"01001011", B"00110100", B"00001101", B"00001101",
 B"00011100", B"11100010", B"00101101", B"00101100", B"00011010",
 B"11101010", B"00011110", B"11011110", B"00100101", B"11101110",
 B"11100010", B"00011100", B"11100001", B"00010010", B"11110100",
 B"00001010", B"00000001", B"11110110", B"11001100", B"00001100",
 B"11011100", B"00011010", B"11011010", B"11111001", B"00101101",
 B"00011000", B"11101000", B"00010111", B"11001001", B"11100000",
 B"11011101", B"00001010", B"00100111", B"00010001", B"00010111",
 B"00100111", B"11000001", B"00010111", B"11001011", B"00000011",
 B"11100110", B"11001001", B"11101001", B"00111010", B"00001010",
 B"00101100", B"00110000", B"11001010", B"11011001", B"11011010",
 B"11000111", B"00000110", B"11011011", B"00101100", B"11111001",
 B"11101010", B"00000110", B"11101010", B"11101011", B"11100100",
 B"00001100", B"00111111", B"11010100", B"01001010", B"11010001",
 B"00011101", B"11101011", B"00111101", B"00011110", B"11110010",
 B"00100001", B"00110101", B"11110000", B"11101111", B"11010010",
 B"00101101", B"11011100", B"00100110", B"11010010", B"11000100",
 B"00100110", B"00010001", B"11000001", B"00011101", B"00100000",
 B"11100011", B"00101000", B"00010011", B"11010010", B"11011101",
 B"00011010", B"11011000", B"11010000", B"11001010", B"00011110",
 B"00101001", B"11001110", B"00100111", B"00011110", B"11110010",
 B"00110000", B"00000111", B"11011000", B"11100010", B"00100001",
 B"11100000", B"11001010", B"11001111", B"00110011", B"00100110",
 B"11011010", B"00001011", B"11010101", B"11100001", B"11110111",
 B"00011011", B"00011110", B"00001001", B"00100010", B"11101111",
 B"11110100", B"00110110", B"11111101", B"11101100", B"00010011",
 B"00001010", B"11100001", B"11010110", B"11110111", B"11011000",
 B"11111111", B"00101000", B"11011110", B"00100011", B"11100000",
 B"11010010", B"00010110", B"00010011", B"00101110", B"00101001",
 B"11110111", B"00010110", B"11011010", B"00011011", B"11101110",
 B"00011110", B"11110101", B"11100011", B"11001110", B"11011000",
 B"00101111", B"11100000", B"00110100", B"00001011", B"00011010",
 B"00010110", B"11110010", B"00111101", B"11100101", B"00101001",
 B"11011111", B"00110000", B"11100101", B"00110011", B"00101100",
 B"11010000", B"00010111", B"00100101", B"11010000", B"00100110",
 B"11100111", B"11101010", B"00100011", B"11101101", B"11010111",
 B"11110101", B"11101101", B"00011101", B"11011000", B"00110001",
 B"00011100", B"11011010", B"00100011", B"00010110", B"11101110",
 B"00100010", B"11001011", B"11110010", B"00101001", B"11011001",
 B"11010110", B"11010100", B"11011100", B"11011001", B"11101110",
 B"11100110", B"00100100", B"00101111", B"11111010", B"00011001",
 B"11101001", B"11010000", B"00110101", B"11010100", B"11000110",
 B"11100100", B"00010011", B"00001001", B"11101110", B"11011000",
 B"00100100", B"11010001", B"00010000", B"11010010", B"11011100",
 B"00010111", B"00010001", B"00100111", B"11010100", B"00001110",
 B"00001001", B"11000111", B"00011001", B"00010100", B"11011100",
 B"11011010", B"00101011", B"11101110", B"11010011", B"11101110",
 B"00110000", B"00111001", B"11011110", B"00011100", B"11011000",
 B"00000111", B"00011101", B"11011000", B"10111010", B"11011010",
 B"11101101", B"11110011", B"00010111", B"11000011", B"00011110",
 B"11010100", B"00000110", B"00011010", B"00101110", B"00111111",
 B"00011000", B"11010111", B"00010011", B"00011010", B"11011110",
 B"11110011", B"00010010", B"11011011", B"11101111", B"00010110",
 B"00111000", B"00010111", B"00011010", B"11100110", B"11101001",
 B"11110111", B"11100001", B"11011100", B"00100010", B"00100011",
 B"11101111", B"00101101", B"11001010", B"00000000", B"00100001",
 B"11100100", B"11101110", B"11111001", B"00011010", B"11101010",
 B"11001100", B"00100000", B"00011010", B"11101101", B"00011100",
 B"00010110", B"11010110", B"11001110", B"00101000", B"00000000",
 B"11000110", B"00110101", B"00011110", B"00010111", B"00100000",
 B"11110001", B"11011011", B"00101000", B"11100100", B"00000111",
 B"00100001", B"11101111", B"11011011", B"11001001", B"11100010",
 B"00101100", B"00100000", B"11011011", B"11100010", B"00100000",
 B"00001000", B"11010011", B"11010100", B"11101100", B"11101100",
 B"11101010", B"00110010", B"00101100", B"11100110", B"00011111",
 B"11100111", B"11100010", B"00110010", B"11100010", B"00011010",
 B"11011101", B"11010111", B"00011011", B"00100011", B"00000011",
 B"11100011", B"00000110", B"11100001", B"11001101", B"00110111",
 B"11001110", B"00100011", B"00110001", B"11011001", B"11110000",
 B"11101111", B"11011110", B"00001010", B"11111000", B"00100110",
 B"00010110", B"00011001", B"11010101", B"00110100", B"00101000",
 B"11101101", B"11100010", B"11111111", B"11001101", B"11100100",
 B"00100011", B"11011100", B"00001110", B"11011111", B"11011011",
 B"00001110", B"11011101", B"01000000", B"00010100", B"00001001",
 B"11110001", B"00001111", B"11110011", B"00101111", B"11011010",
 B"11111001", B"11001010", B"11011110", B"00111111", B"00000000",
 B"00111010", B"00100101", B"11001111", B"00011000", B"11101000",
 B"00011010", B"11001001", B"11110111", B"00011100", B"00011000",
 B"11010100", B"11110100", B"00011110", B"11000110", B"00100110",
 B"11010000", B"11011101", B"00011101", B"11010111", B"00110100",
 B"01000000", B"11110100", B"11100000", B"11011111", B"11100110",
 B"11100110", B"11100111", B"00011100", B"00110001", B"11100010",
 B"00100011", B"11100010", B"11100000", B"11111111", B"00100111",
 B"11100000", B"11100100", B"00010010", B"11001001", B"11000010",
 B"11100110", B"11100101", B"11101001", B"00011001", B"11011111",
 B"00101110", B"11001100", B"11101011", B"00010001", B"11111001",
 B"00101111", B"00011011", B"11011100", B"11010011", B"00001001",
 B"00100011", B"11100000", B"11110000", B"00011111", B"00011001",
 B"11100001", B"00000100", B"00100111", B"11101101", B"11100100",
 B"00011101", B"11010010", B"00100001", B"00011000", B"11010100",
 B"11011001", B"11011100", B"11100010", B"11100011", B"00011111",
 B"00010011", B"00001110", B"00011110", B"00100011", B"00011011",
 B"00010100", B"00110000", B"00101000", B"11001101", B"00100000",
 B"11111010", B"11100111", B"11100101", B"00011101", B"00110101",
 B"11111110", B"11010101", B"00011101", B"00011010", B"11101011",
 B"00100110", B"00010001", B"11101101", B"10111110", B"00010110",
 B"11010101", B"00101100", B"11100100", B"11010010", B"00000110",
 B"00001100", B"11101100", B"11011110", B"11110001", B"00101001",
 B"00110100", B"11001100", B"00100010", B"11101000", B"11011101",
 B"00101101", B"00001001", B"00000101", B"11110010", B"11100000",
 B"11100011", B"11011001", B"00010000", B"11100011", B"11001010",
 B"00010011", B"11011000", B"11101011", B"11011111", B"11101110",
 B"11001111", B"00011001", B"11001100", B"11110111", B"11100010",
 B"00110010", B"00001100", B"11011111", B"11100011", B"00111100",
 B"00100010", B"00011001", B"11101001", B"00100110", B"11100110",
 B"00110011", B"11011101", B"11000010", B"00111010", B"11100000",
 B"00100110", B"11111011", B"11100111", B"00010101", B"11010100",
 B"00011100", B"11011010", B"00101111", B"11011101", B"11011001",
 B"00110101", B"11111110", B"00011111", B"00100000", B"11101011",
 B"00101111", B"00011000", B"11001110", B"11011000", B"00101011",
 B"11010010", B"11101111", B"11011001", B"11010110", B"00011001",
 B"00011110", B"00010101", B"00110110", B"11010110", B"00101001",
 B"00110010", B"00011100", B"11100010", B"00100111", B"11010100",
 B"00100111", B"11110010", B"00100110", B"11010011", B"11001100",
 B"11100101", B"00110100", B"00100011", B"11100011", B"00001111",
 B"11000101", B"11001000", B"00101001", B"11100010", B"11011001",
 B"11010101", B"11011000", B"11111101", B"00111000", B"00100011",
 B"00100101", B"11110111", B"00100101", B"11011101", B"00110001",
 B"11011110", B"00001011", B"11011100", B"00001110", B"11011100",
 B"11011101", B"00110001", B"00101000", B"00110111", B"00001000",
 B"11010111", B"00011100", B"00011011", B"11100010", B"11011000",
 B"00110100", B"11011010", B"11011001", B"00100001", B"00010111",
 B"00111001", B"00101111", B"11001110", B"11000100", B"00010101",
 B"00101010", B"00011000", B"00001111", B"00011011", B"00010110",
 B"00100110", B"01000000", B"11100101", B"00011100", B"00100101",
 B"11011111", B"11011000", B"11101111", B"11101010", B"11100001",
 B"00101001", B"11011100", B"11011101", B"00100101", B"11010100",
 B"11010011", B"11011111", B"11011111", B"11101011", B"11100001",
 B"11011001", B"11110111", B"00010111", B"00100011", B"00110010",
 B"00011100", B"11001110", B"00001111", B"00110000", B"00101001",
 B"11011000", B"00101100", B"11011100", B"00010011", B"00110110",
 B"11010111", B"00101101", B"00011110", B"11010010", B"00001101",
 B"00010100", B"11000011", B"11100100", B"11100000", B"11001011",
 B"11111100", B"00110100", B"00101000", B"00100000", B"00001001",
 B"11110110", B"11110101", B"11110001", B"11011011", B"00101101",
 B"11011100", B"10111011", B"00001001", B"11101100", B"00101110",
 B"11001001", B"11011011", B"10111110", B"00011101", B"00110010",
 B"11101111", B"00001101", B"11110111", B"00001011", B"00011010",
 B"00100111", B"00010101", B"00010001", B"00001100", B"11011000",
 B"00011000", B"11000000", B"00001101", B"11111110", B"11100000",
 B"00110011", B"00111000", B"00100001", B"00110001", B"00110011",
 B"11101000", B"00100000", B"11011011", B"00100100", B"11100111",
 B"00101001", B"00010110", B"11001010", B"11010110", B"00000011",
 B"00010110", B"11011101", B"11011100", B"00000011", B"00100010",
 B"11100100", B"11100010", B"11101000", B"11101110", B"01000100",
 B"11100110", B"11101110", B"00011000", B"11100011", B"00000000",
 B"11010100", B"00001111", B"00011110", B"11010010", B"00111100",
 B"00011100", B"11011011", B"00011100", B"00011101", B"11011101",
 B"11101001", B"00100010", B"00101000", B"11100110", B"11001001",
 B"11110000", B"11010101", B"11110010", B"11110001", B"11100111",
 B"11011010", B"00011111", B"11011000", B"00011011", B"11011001",
 B"11110110", B"00001100", B"00011111", B"11011111", B"11111100",
 B"00010001", B"00100001", B"11101011", B"00011110", B"11010101",
 B"00011110", B"11100110", B"11011100", B"11010011", B"00101000",
 B"00100111", B"11011110", B"00110010", B"11100110", B"00100110",
 B"11110000", B"00101101", B"11110011", B"11100000", B"11101011",
 B"00110100", B"00011110", B"11101100", B"00101000", B"11101010",
 B"11111110", B"11001111", B"11100011", B"00101101", B"00100001",
 B"11100110", B"11010101", B"00100011", B"00100110", B"00111101",
 B"00100111", B"11100111", B"11011001", B"11010111", B"00011011",
 B"10111101", B"00111011", B"11100011", B"11001001", B"01000101",
 B"00000101", B"11011100", B"11101010", B"10110001", B"00001001",
 B"00011101", B"11011011", B"00110101", B"11101110", B"11010011",
 B"11010001", B"00011011", B"11011000", B"00100001", B"11100010",
 B"11100100", B"00011111", B"00100110", B"00101100", B"00001111",
 B"11000100", B"11110001", B"11100000", B"00110000", B"11011110",
 B"00000100", B"11100111", B"00011111", B"11001010", B"11010011",
 B"11011101", B"00100101", B"00010011", B"00011101", B"00100110",
 B"00001001", B"11010110", B"00101000", B"11011011", B"00001100",
 B"11110001", B"00101111", B"11110010", B"11100011", B"00011000",
 B"11111001", B"11000011", B"11100110", B"11110101", B"11100101",
 B"11011001", B"00001111", B"11010111", B"00111001", B"11100101",
 B"10111010", B"00101110", B"11111111", B"11100000", B"11101101",
 B"11100001", B"11110001", B"00001100", B"11101101", B"00101110",
 B"11011110", B"11010111", B"00011001", B"00010011", B"00100000",
 B"00100111", B"11100110", B"11100100", B"11101011", B"11100110",
 B"11110001", B"11100001", B"00001110", B"00101010", B"01000000",
 B"00110000", B"11011001", B"11011000", B"11101011", B"11000011",
 B"11111111", B"00111000", B"00100000", B"00011001", B"00100001",
 B"00101010", B"11100111", B"11011111", B"11111110", B"00100101",
 B"11001010", B"11000011", B"00000010", B"11001111", B"11111100",
 B"11010010", B"11100100", B"00101101", B"11000010", B"00100010",
 B"00100010", B"00001010", B"00101110", B"00110101", B"00000100",
 B"00000101", B"00011101", B"00100011", B"00110000", B"11010111",
 B"11011000", B"00101111", B"11011001", B"11111110", B"11101010",
 B"11100100", B"00100011", B"11011110", B"00101110", B"00010101",
 B"11000100", B"00001110", B"00100111", B"11110101", B"11001010",
 B"00010101", B"00000111", B"11001100", B"11011010", B"11101111",
 B"11000010", B"11101110", B"11101000", B"00001110", B"00001101",
 B"11100000", B"11011011", B"11001110", B"11101000", B"11010011",
 B"00111110", B"11001111", B"00011101", B"00011010", B"11100000",
 B"00011111", B"00100111", B"11011111", B"00011111", B"00001011",
 B"11110011", B"01001001", B"00101001", B"11000111", B"11110101",
 B"00100011", B"10111111", B"00101100", B"11001101", B"11100101",
 B"11001110", B"00001101", B"00000001", B"00001001", B"00101010",
 B"01000101", B"11000010", B"00101010", B"00100000", B"11100111",
 B"11100111", B"00001010", B"11101000", B"11101101", B"00011000",
 B"11110010", B"00010011", B"11001001", B"11101001", B"00010110",
 B"01000100", B"00010110", B"00100100", B"01000011", B"00010010",
 B"00010100", B"00011101", B"00101001", B"11111110", B"11111111",
 B"11101110", B"00001010", B"00001101", B"11100010", B"00101111",
 B"11101111", B"00010001", B"11100010", B"11111010", B"00101001",
 B"11101001", B"00001101", B"11001101", B"11111000", B"11101010",
 B"11010011", B"11011011", B"11010000", B"00110110", B"01000000",
 B"00001101", B"00100011", B"11101000", B"11000111", B"00011100",
 B"11011110", B"00101001", B"11010010", B"11001111", B"00101111",
 B"00100000", B"00001110", B"11010010", B"11101010", B"00010000",
 B"00001101", B"11001111", B"11010010", B"00010110", B"11011111",
 B"11100100", B"11011010", B"11000100", B"00101110", B"10111101",
 B"00000010", B"11001011", B"11110010", B"00100010", B"00011101",
 B"00101101", B"00111011", B"11100110", B"11101101", B"11100011",
 B"11100001", B"11101111", B"00001100", B"00111000", B"11100000",
 B"00100111", B"11111001", B"11011111", B"00011011", B"11101100",
 B"11100100", B"11000101", B"00001010", B"00011101", B"11110001",
 B"11101000", B"11011010", B"00010100", B"11100011", B"00100111",
 B"11001000", B"11101001", B"00010010", B"00100110", B"00101000",
 B"00011011", B"11010111", B"00101010", B"11011111", B"00011011",
 B"11001001", B"10111000", B"11011001", B"00010101", B"11110110",
 B"00101100", B"11011000", B"11100001", B"00001111", B"00110000",
 B"00101111", B"11011110", B"11010011", B"00100000", B"00101000",
 B"11010101", B"11100001", B"00100010", B"00011110", B"11000011",
 B"00110000", B"11111010", B"11101100", B"11101101", B"00100101",
 B"11011110", B"00001011", B"11101101", B"11011110", B"11111001",
 B"00010111", B"00110000", B"11001111", B"00100000", B"00011100",
 B"11111101", B"11011101", B"00001100", B"00100011", B"11010100",
 B"11010010", B"00101011", B"00101110", B"00111011", B"11000100",
 B"00110100", B"11101001", B"00100011", B"11101110", B"11101011",
 B"11001100", B"00100011", B"00000001", B"00011001", B"00010011",
 B"11101001", B"11001010", B"00100011", B"00001110", B"00100000",
 B"11011000", B"00011101", B"11011100", B"00100111", B"11011110",
 B"11100110", B"00100010", B"11010011", B"11100010", B"11001110",
 B"00011010", B"00100110", B"11001001", B"00100011", B"11111110",
 B"11011111", B"11010011", B"11100011", B"00100001", B"11100101",
 B"00100000", B"00011001", B"11011111", B"00101111", B"11110000",
 B"11100010", B"11011111", B"00101001", B"00100010", B"11001010",
 B"00011110", B"11011111", B"00010111", B"11001011", B"11001000",
 B"00011101", B"00010001", B"00000000", B"00110010", B"11010110",
 B"00001000", B"10111111", B"11110110", B"00101101", B"00010110",
 B"00011011", B"00101001", B"00100100", B"11100000", B"00110100",
 B"11101111", B"00101001", B"11110000", B"00101110", B"00011101",
 B"11010100", B"10110101", B"00010001", B"00100001", B"11011110",
 B"11001000", B"11011100", B"11100101", B"11100011", B"00100011",
 B"00101001", B"11101011", B"00100101", B"11000111", B"00110110",
 B"00110110", B"00011101", B"11111111", B"00111011", B"00100011",
 B"00110101", B"00010000", B"11010000", B"11011110", B"00110010",
 B"00101000", B"00100011", B"00100000", B"11101100", B"11110011",
 B"00101100", B"11011010", B"00001000", B"11001000", B"11011111",
 B"00100011", B"11110010", B"00100011", B"00010110", B"00010110",
 B"00111100", B"11011111", B"00101101", B"11101100", B"00010111",
 B"11011111", B"11110100", B"00110011", B"00011100", B"00101001",
 B"11101101", B"00011100", B"11100001", B"00101010", B"00011010",
 B"00011101", B"11101010", B"00110111", B"00010111", B"00000011",
 B"11011110", B"00100001", B"01010011", B"00011000", B"00101000",
 B"00100111", B"00100101", B"00100010", B"00011100", B"00101001",
 B"11101001", B"11010110", B"11100100", B"10111110", B"00110011",
 B"00011000", B"00101001", B"00011101", B"00110100", B"00101011",
 B"11101010", B"00101001", B"00111000", B"11100001", B"11011110",
 B"00100110", B"11110100", B"11101000", B"11011100", B"00100110",
 B"00101010", B"11001000", B"00001011", B"11011101", B"00100010",
 B"11011000", B"11100010", B"11011111", B"11101100", B"00011000",
 B"11100001", B"00010001", B"11111101", B"11010001", B"00110101",
 B"11110010", B"00110001", B"11110011", B"11100000", B"00101011",
 B"00101010", B"00110110", B"11011011", B"11110010", B"00100010",
 B"00110010", B"10111100", B"11101100", B"11111010", B"11101010",
 B"00011110", B"11110001", B"00001111", B"11100100", B"11011111",
 B"00001110", B"11000001", B"00100000", B"00010101", B"11110100",
 B"11110011", B"11010011", B"11101101", B"11001101", B"00110010",
 B"00011110", B"00100001", B"10111101", B"00100110", B"11011111",
 B"00110100", B"11110101", B"00111011", B"11111010", B"11101000",
 B"11001100", B"11100110", B"00001111", B"11101001", B"00010010",
 B"11010100", B"00101001", B"11011100", B"11000101", B"11011101",
 B"00100001", B"00011111", B"11100000", B"00101110", B"11110111",
 B"00011100", B"11110100", B"11101000", B"11110010", B"00001010",
 B"00111000", B"00101001", B"11101100", B"11100001", B"11001111",
 B"00001000", B"00011000", B"11101001", B"00010000", B"00100010",
 B"00010111", B"11011111", B"00010101", B"00010110", B"10111010",
 B"11101101", B"00001000", B"00100101", B"11100010", B"00010101",
 B"00011000", B"11101001", B"00010100", B"00010010", B"11011100",
 B"00101110", B"00111000", B"11100001", B"11110100", B"00100000",
 B"00000101", B"11010010", B"11011110", B"11100000", B"00011010",
 B"11001000", B"11011011", B"11101011", B"00100110", B"00011100",
 B"11100000", B"11001111", B"11011001", B"00000000", B"00100000",
 B"00101010", B"11101000", B"00001100", B"11110011", B"11001000",
 B"11000101", B"11011110", B"00101110", B"00010000", B"11101010",
 B"00101100", B"11100110", B"11100001", B"11010001", B"11110011",
 B"00001101", B"00011000", B"00010100", B"00010000", B"00001100",
 B"11101111", B"11110000", B"00110011", B"11101101", B"00110000",
 B"11100011", B"11010000", B"00100101", B"11010111", B"11001100",
 B"11100101", B"00101000", B"00000111", B"11010110", B"00101010",
 B"11100100", B"11101100", B"00010000", B"00101010", B"11010010",
 B"11001011", B"11100110", B"11001100", B"11011000", B"11100010",
 B"00011101", B"11100110", B"11111001", B"11000101", B"00100101",
 B"00100111", B"11011001", B"00011000", B"11000101", B"11111001",
 B"00010011", B"11101110", B"00110100", B"00100111", B"11110001",
 B"00111010", B"00011000", B"11100000", B"11011000", B"00001101",
 B"00000100", B"11100111", B"11111100", B"11110000", B"00010101",
 B"00001101", B"11010101", B"11100010", B"10111011", B"11011110",
 B"11100100", B"00101110", B"00101000", B"11101101", B"11011110",
 B"00100101", B"00001111", B"11111010", B"11011110", B"11110011",
 B"11110011", B"11010010", B"11110001", B"00110100", B"00011001",
 B"00011110", B"00011100", B"00001100", B"11001111", B"00010101",
 B"00010101", B"11011110", B"00100111", B"00100101", B"11100100",
 B"11101011", B"00011101", B"00011001", B"00101000", B"11100000",
 B"00100000", B"11101010", B"00001110", B"11010101", B"11101101",
 B"11011100", B"00110000", B"11111101", B"11100101", B"00011110",
 B"11011000", B"11011100", B"01000101", B"00100110", B"11010011",
 B"11100110", B"11100011", B"11110110", B"11110010", B"11101111",
 B"11000000", B"11011101", B"11011101", B"00110110", B"00110010",
 B"00101010", B"00100100", B"11001000", B"11110110", B"11011111",
 B"00100010", B"00100101", B"11011010", B"00110101", B"11100101",
 B"11010011", B"11010010", B"00110000", B"00100001", B"00011101",
 B"00001101", B"11100000", B"11011101", B"11100011", B"00011101",
 B"11010001", B"11001011", B"11100110", B"00100100", B"00011010",
 B"11111000", B"00010110", B"11010101", B"11011001", B"11011101",
 B"11101100", B"00100110", B"11011100", B"00110110", B"11010001",
 B"00100100", B"00010010", B"11011010", B"11101111", B"11010101",
 B"11111001", B"11101111", B"00011000", B"00110101", B"00101101",
 B"00110110", B"00010101", B"00011110", B"00001111", B"00101010",
 B"00010100", B"11010110", B"00011110", B"00101001", B"11110001",
 B"00001111", B"00010000", B"11011001", B"11101011", B"00001111",
 B"11011000", B"00100000", B"11110001", B"11100101", B"00100111",
 B"00100010", B"00100100", B"11100010", B"00001001", B"11011000",
 B"11011111", B"11111101", B"00101111", B"00100110", B"00111100",
 B"00010110", B"11100100", B"00101101", B"00000010", B"11100101",
 B"11011000", B"11101110", B"11100000", B"00000101", B"00100001",
 B"11010001", B"11100111", B"11010001", B"11110000", B"11011011",
 B"00011111", B"11011111", B"11011010", B"00100001", B"11110100",
 B"11111110", B"11001101", B"11100100", B"00010110", B"11011000",
 B"11001000", B"11100001", B"11001001", B"00011010", B"11101010",
 B"00100101", B"11101100", B"11101001", B"11110001", B"11010100",
 B"00010111", B"00110100", B"00000110", B"00110001", B"00001111",
 B"10111011", B"11011001", B"11101111", B"11110001", B"00101100",
 B"11100111", B"00011000", B"00101110", B"11011110", B"11011010",
 B"00011101", B"11001110", B"11011000", B"11001101", B"00001100",
 B"11011111", B"00110110", B"01000011", B"00011111", B"11010000",
 B"00010111", B"11101111", B"00101111", B"11110100", B"11011000",
 B"00100110", B"11011101", B"00100000", B"11001100", B"11011001",
 B"00011011", B"00110011", B"00010001", B"11010001", B"11100000",
 B"00101011", B"00011111", B"11001110", B"11100000", B"00101000",
 B"11101010", B"11110000", B"11010100", B"11010101", B"00010011",
 B"11100010", B"00101001", B"11001100", B"11110011", B"00101010",
 B"11110100", B"00100000", B"11010000", B"11110001", B"00011000",
 B"11100000", B"00101010", B"11110111", B"11110100", B"11110111",
 B"00010001", B"00000010", B"11001001", B"00000110", B"00111001",
 B"00100111", B"00100000", B"00101111", B"00101110", B"00101100",
 B"00010111", B"00100011", B"00101101", B"00011000", B"00011001",
 B"00100011", B"00100010", B"00000000", B"00011111", B"11000011",
 B"11110110", B"00011111", B"11100101", B"00101110", B"11011011",
 B"11100000", B"00001110", B"00011110", B"11001101", B"00011111",
 B"00100000", B"11011011", B"00011010", B"00011110", B"11100110",
 B"11010110", B"11010001", B"11100111", B"00000111", B"00101101",
 B"11101110", B"00100110", B"11010011", B"11111111", B"11100000",
 B"11010111", B"00101001", B"11011010", B"11101110", B"11010010",
 B"11100001", B"11100000", B"00011000", B"11100101", B"00101011",
 B"11010001", B"11101010", B"00010101", B"00001110", B"11110110",
 B"11101111", B"00100011", B"00110111", B"11100011", B"00101001",
 B"00011110", B"11001110", B"11011101", B"10110011", B"00000010",
 B"11111000", B"00011110", B"00100111", B"00101000", B"00101001",
 B"11001111", B"00000110", B"11001110", B"00010111", B"11001011",
 B"11101010", B"00100011", B"00101001", B"11010010", B"11011000",
 B"00011010", B"11001111", B"00100000", B"11001010", B"11010001",
 B"00011011", B"11100010", B"11100001", B"00001000", B"11101101",
 B"00011111", B"11011011", B"11100101", B"00001101", B"00011001",
 B"11100000", B"11100100", B"01000101", B"11011001", B"11101010",
 B"11001001", B"11100110", B"11010111", B"11101001", B"00011010",
 B"00101001", B"00011111", B"00111101", B"11110000", B"11001000"

);

signal input_counter : integer range 0 to 19999 := 0;
signal start_fifo    : bit_vector (7 downto 0) := ( B"0100_0000" );
signal clk : bit;

begin

process (clk, clear)
begin
if (clear = '1') then
    rxin <= (others => '0');
elsif (clk = '1' and clk'event) then
    rxin <= input_bank(input_counter);
end if;
end process;

process (clk, clear)
begin
if (clear = '1') then
    input_counter <= 0;
elsif (clk = '1' and clk'event) then
    if (input_counter < 19999) then
    input_counter <= input_counter + 1;
    else
    input_counter <= 0;
    end if;
end if;
end process;

rom_pos <= input_counter;

process (clk, clear)
begin
if (clear = '1') then
    start_fifo <= B"0100_0000";
elsif ( clk = '1' and clk'event) then
    start_fifo <= start_fifo (6 downto 0) & start_fifo (7);
end if;
end process;

clk   <= clock;
start <= start_fifo (7);

end test_bench;
